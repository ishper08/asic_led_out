magic
tech sky130A
magscale 1 2
timestamp 1680496449
<< obsli1 >>
rect 1104 2159 18860 47345
<< obsm1 >>
rect 750 2128 19019 47376
<< metal2 >>
rect 4986 0 5042 800
rect 14922 0 14978 800
<< obsm2 >>
rect 756 856 19013 47977
rect 756 800 4930 856
rect 5098 800 14866 856
rect 15034 800 19013 856
<< metal3 >>
rect 0 47880 800 48000
rect 0 44344 800 44464
rect 0 40808 800 40928
rect 0 37272 800 37392
rect 0 33736 800 33856
rect 0 30200 800 30320
rect 0 26664 800 26784
rect 0 23128 800 23248
rect 0 19592 800 19712
rect 0 16056 800 16176
rect 0 12520 800 12640
rect 0 8984 800 9104
rect 0 5448 800 5568
rect 0 1912 800 2032
<< obsm3 >>
rect 880 47800 19017 47973
rect 800 44544 19017 47800
rect 880 44264 19017 44544
rect 800 41008 19017 44264
rect 880 40728 19017 41008
rect 800 37472 19017 40728
rect 880 37192 19017 37472
rect 800 33936 19017 37192
rect 880 33656 19017 33936
rect 800 30400 19017 33656
rect 880 30120 19017 30400
rect 800 26864 19017 30120
rect 880 26584 19017 26864
rect 800 23328 19017 26584
rect 880 23048 19017 23328
rect 800 19792 19017 23048
rect 880 19512 19017 19792
rect 800 16256 19017 19512
rect 880 15976 19017 16256
rect 800 12720 19017 15976
rect 880 12440 19017 12720
rect 800 9184 19017 12440
rect 880 8904 19017 9184
rect 800 5648 19017 8904
rect 880 5368 19017 5648
rect 800 2112 19017 5368
rect 880 1939 19017 2112
<< metal4 >>
rect 3163 2128 3483 47376
rect 5382 2128 5702 47376
rect 7602 2128 7922 47376
rect 9821 2128 10141 47376
rect 12041 2128 12361 47376
rect 14260 2128 14580 47376
rect 16480 2128 16800 47376
rect 18699 2128 19019 47376
<< obsm4 >>
rect 1899 5475 3083 30429
rect 3563 5475 5302 30429
rect 5782 5475 7522 30429
rect 8002 5475 8221 30429
<< labels >>
rlabel metal2 s 4986 0 5042 800 6 clk
port 1 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 led_out[0]
port 2 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 led_out[1]
port 3 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 led_out[2]
port 4 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 led_out[3]
port 5 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 led_out[4]
port 6 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 led_out[5]
port 7 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 led_out[6]
port 8 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 led_out_b[0]
port 9 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 led_out_b[1]
port 10 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 led_out_b[2]
port 11 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 led_out_b[3]
port 12 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 led_out_b[4]
port 13 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 led_out_b[5]
port 14 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 led_out_b[6]
port 15 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 reset
port 16 nsew signal input
rlabel metal4 s 3163 2128 3483 47376 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 47376 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 47376 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 47376 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 47376 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 47376 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 47376 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 47376 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1333090
string GDS_FILE /home/ish/work/caravel/caravel_walkthrough/openlane/segment7/runs/23_04_03_14_31/results/signoff/segment7.magic.gds
string GDS_START 435278
<< end >>

