magic
tech sky130A
magscale 1 2
timestamp 1680496446
<< viali >>
rect 1593 47141 1627 47175
rect 1777 46937 1811 46971
rect 1593 44829 1627 44863
rect 1777 41089 1811 41123
rect 1593 40953 1627 40987
rect 1593 37621 1627 37655
rect 6837 36193 6871 36227
rect 6377 36125 6411 36159
rect 6745 36125 6779 36159
rect 5917 36057 5951 36091
rect 4629 35649 4663 35683
rect 4813 35649 4847 35683
rect 4721 35445 4755 35479
rect 6101 35037 6135 35071
rect 6929 35037 6963 35071
rect 6377 34901 6411 34935
rect 6561 34561 6595 34595
rect 7297 34561 7331 34595
rect 7481 34561 7515 34595
rect 6745 34357 6779 34391
rect 6285 34153 6319 34187
rect 7573 34153 7607 34187
rect 6837 34085 6871 34119
rect 6193 34017 6227 34051
rect 6655 33949 6689 33983
rect 1593 33881 1627 33915
rect 1777 33881 1811 33915
rect 7557 33881 7591 33915
rect 7757 33881 7791 33915
rect 6653 33813 6687 33847
rect 7389 33813 7423 33847
rect 7297 33065 7331 33099
rect 5457 32997 5491 33031
rect 7481 32929 7515 32963
rect 5733 32861 5767 32895
rect 6377 32861 6411 32895
rect 7573 32861 7607 32895
rect 7941 32725 7975 32759
rect 5181 32385 5215 32419
rect 5365 32385 5399 32419
rect 5457 32385 5491 32419
rect 5549 32385 5583 32419
rect 5825 32181 5859 32215
rect 5273 31773 5307 31807
rect 5917 31773 5951 31807
rect 5917 31433 5951 31467
rect 5457 31297 5491 31331
rect 6009 31297 6043 31331
rect 6745 31297 6779 31331
rect 6837 31297 6871 31331
rect 7021 31297 7055 31331
rect 7113 31297 7147 31331
rect 6561 31093 6595 31127
rect 1593 30685 1627 30719
rect 6009 30685 6043 30719
rect 6101 30685 6135 30719
rect 6469 30685 6503 30719
rect 7113 30685 7147 30719
rect 7481 30685 7515 30719
rect 8033 30685 8067 30719
rect 5733 30617 5767 30651
rect 8217 30549 8251 30583
rect 7021 30209 7055 30243
rect 7297 30209 7331 30243
rect 7481 30209 7515 30243
rect 8033 30209 8067 30243
rect 7389 30073 7423 30107
rect 8125 30005 8159 30039
rect 5641 29801 5675 29835
rect 7481 29801 7515 29835
rect 4905 29597 4939 29631
rect 6193 29597 6227 29631
rect 6745 29597 6779 29631
rect 6929 29597 6963 29631
rect 7573 29597 7607 29631
rect 5181 29529 5215 29563
rect 4629 29461 4663 29495
rect 4813 29461 4847 29495
rect 4997 29461 5031 29495
rect 7941 29257 7975 29291
rect 5181 29121 5215 29155
rect 6561 29121 6595 29155
rect 6653 29121 6687 29155
rect 6837 29121 6871 29155
rect 6929 29121 6963 29155
rect 7757 29121 7791 29155
rect 8033 29121 8067 29155
rect 4905 29053 4939 29087
rect 4997 29053 5031 29087
rect 5089 29053 5123 29087
rect 7573 28985 7607 29019
rect 4721 28917 4755 28951
rect 7113 28917 7147 28951
rect 4445 28713 4479 28747
rect 4813 28645 4847 28679
rect 6469 28577 6503 28611
rect 6653 28577 6687 28611
rect 8033 28577 8067 28611
rect 3249 28509 3283 28543
rect 3433 28509 3467 28543
rect 6561 28509 6595 28543
rect 6745 28509 6779 28543
rect 7481 28509 7515 28543
rect 7665 28509 7699 28543
rect 4445 28441 4479 28475
rect 3341 28373 3375 28407
rect 4261 28373 4295 28407
rect 6285 28373 6319 28407
rect 7941 28373 7975 28407
rect 8585 28033 8619 28067
rect 8861 28033 8895 28067
rect 8493 27965 8527 27999
rect 3341 27557 3375 27591
rect 3433 27489 3467 27523
rect 3157 27421 3191 27455
rect 3249 27421 3283 27455
rect 3985 27421 4019 27455
rect 4261 27421 4295 27455
rect 4445 27421 4479 27455
rect 4629 27421 4663 27455
rect 4813 27353 4847 27387
rect 4629 27081 4663 27115
rect 6561 27013 6595 27047
rect 6929 27013 6963 27047
rect 7021 27013 7055 27047
rect 1777 26945 1811 26979
rect 4445 26945 4479 26979
rect 5641 26945 5675 26979
rect 5733 26945 5767 26979
rect 7113 26945 7147 26979
rect 4261 26877 4295 26911
rect 7297 26877 7331 26911
rect 8033 26877 8067 26911
rect 1593 26809 1627 26843
rect 8309 26809 8343 26843
rect 5917 26741 5951 26775
rect 8493 26741 8527 26775
rect 4353 26537 4387 26571
rect 4537 26537 4571 26571
rect 6653 26469 6687 26503
rect 4997 26401 5031 26435
rect 7021 26401 7055 26435
rect 4537 26333 4571 26367
rect 4905 26333 4939 26367
rect 5825 26333 5859 26367
rect 6009 26333 6043 26367
rect 6837 26333 6871 26367
rect 6929 26333 6963 26367
rect 7113 26333 7147 26367
rect 6193 26265 6227 26299
rect 6561 25993 6595 26027
rect 3985 25857 4019 25891
rect 4169 25857 4203 25891
rect 6745 25857 6779 25891
rect 6837 25789 6871 25823
rect 6929 25789 6963 25823
rect 7021 25789 7055 25823
rect 4169 25653 4203 25687
rect 2145 25449 2179 25483
rect 6285 25449 6319 25483
rect 6469 25449 6503 25483
rect 8125 25449 8159 25483
rect 5549 25313 5583 25347
rect 5365 25245 5399 25279
rect 5825 25245 5859 25279
rect 7849 25245 7883 25279
rect 2329 25177 2363 25211
rect 6437 25177 6471 25211
rect 6653 25177 6687 25211
rect 8309 25177 8343 25211
rect 1961 25109 1995 25143
rect 2145 25109 2179 25143
rect 5733 25109 5767 25143
rect 8125 25109 8159 25143
rect 3893 24905 3927 24939
rect 5273 24905 5307 24939
rect 7925 24837 7959 24871
rect 8125 24837 8159 24871
rect 5181 24769 5215 24803
rect 5457 24769 5491 24803
rect 6745 24769 6779 24803
rect 7021 24769 7055 24803
rect 3525 24701 3559 24735
rect 6837 24701 6871 24735
rect 4077 24633 4111 24667
rect 6561 24633 6595 24667
rect 7757 24633 7791 24667
rect 3893 24565 3927 24599
rect 7021 24565 7055 24599
rect 7941 24565 7975 24599
rect 4169 24361 4203 24395
rect 5641 24361 5675 24395
rect 8033 24293 8067 24327
rect 4353 24225 4387 24259
rect 4537 24225 4571 24259
rect 1869 24157 1903 24191
rect 2145 24157 2179 24191
rect 4445 24157 4479 24191
rect 4629 24157 4663 24191
rect 5181 24157 5215 24191
rect 5549 24157 5583 24191
rect 5733 24157 5767 24191
rect 6929 24157 6963 24191
rect 7389 24157 7423 24191
rect 7941 24157 7975 24191
rect 8217 24157 8251 24191
rect 7205 24089 7239 24123
rect 1961 24021 1995 24055
rect 2329 24021 2363 24055
rect 5365 24021 5399 24055
rect 8401 24021 8435 24055
rect 7573 23817 7607 23851
rect 4077 23681 4111 23715
rect 4261 23681 4295 23715
rect 7113 23681 7147 23715
rect 7757 23681 7791 23715
rect 7941 23681 7975 23715
rect 6837 23613 6871 23647
rect 4353 23545 4387 23579
rect 1593 23477 1627 23511
rect 5917 23273 5951 23307
rect 6837 23273 6871 23307
rect 5825 23205 5859 23239
rect 5733 23137 5767 23171
rect 6009 23069 6043 23103
rect 6561 23001 6595 23035
rect 5733 22729 5767 22763
rect 5825 22729 5859 22763
rect 7481 22729 7515 22763
rect 8217 22729 8251 22763
rect 5273 22661 5307 22695
rect 5641 22661 5675 22695
rect 1593 22593 1627 22627
rect 1685 22593 1719 22627
rect 6009 22593 6043 22627
rect 7113 22593 7147 22627
rect 7297 22593 7331 22627
rect 8309 22593 8343 22627
rect 8493 22593 8527 22627
rect 1869 22525 1903 22559
rect 1777 22389 1811 22423
rect 4445 22185 4479 22219
rect 5641 21981 5675 22015
rect 7481 21981 7515 22015
rect 7665 21981 7699 22015
rect 4629 21913 4663 21947
rect 5089 21913 5123 21947
rect 5457 21913 5491 21947
rect 5825 21913 5859 21947
rect 7849 21913 7883 21947
rect 4261 21845 4295 21879
rect 4429 21845 4463 21879
rect 5549 21845 5583 21879
rect 5365 21641 5399 21675
rect 5549 21505 5583 21539
rect 5733 21505 5767 21539
rect 5825 21505 5859 21539
rect 7297 21505 7331 21539
rect 7665 21505 7699 21539
rect 8033 21505 8067 21539
rect 8401 21505 8435 21539
rect 8769 21505 8803 21539
rect 7481 21369 7515 21403
rect 2053 21097 2087 21131
rect 5089 21097 5123 21131
rect 8217 21097 8251 21131
rect 1869 20961 1903 20995
rect 2881 20961 2915 20995
rect 2145 20893 2179 20927
rect 3341 20893 3375 20927
rect 5365 20893 5399 20927
rect 8125 20893 8159 20927
rect 3249 20825 3283 20859
rect 5273 20825 5307 20859
rect 5825 20825 5859 20859
rect 1869 20757 1903 20791
rect 3157 20757 3191 20791
rect 5273 20553 5307 20587
rect 5365 20485 5399 20519
rect 3709 20417 3743 20451
rect 5273 20417 5307 20451
rect 5549 20417 5583 20451
rect 3433 20349 3467 20383
rect 3525 20213 3559 20247
rect 3893 20213 3927 20247
rect 2973 20009 3007 20043
rect 2605 19941 2639 19975
rect 1777 19805 1811 19839
rect 1593 19737 1627 19771
rect 2973 19737 3007 19771
rect 3157 19669 3191 19703
rect 2795 19465 2829 19499
rect 2697 19397 2731 19431
rect 2881 19397 2915 19431
rect 1777 19329 1811 19363
rect 2053 19329 2087 19363
rect 2145 19329 2179 19363
rect 2973 19329 3007 19363
rect 1593 19261 1627 19295
rect 3157 18921 3191 18955
rect 3341 18921 3375 18955
rect 5917 18921 5951 18955
rect 2973 18785 3007 18819
rect 3157 18717 3191 18751
rect 4997 18717 5031 18751
rect 5365 18717 5399 18751
rect 2881 18649 2915 18683
rect 2053 18241 2087 18275
rect 2881 18241 2915 18275
rect 2973 18241 3007 18275
rect 2237 18173 2271 18207
rect 2789 18173 2823 18207
rect 3065 18173 3099 18207
rect 1869 18037 1903 18071
rect 3249 18037 3283 18071
rect 2973 17833 3007 17867
rect 3341 17833 3375 17867
rect 2145 17697 2179 17731
rect 3065 17697 3099 17731
rect 2329 17629 2363 17663
rect 2421 17629 2455 17663
rect 3157 17629 3191 17663
rect 2881 17561 2915 17595
rect 2145 17493 2179 17527
rect 2881 17153 2915 17187
rect 3065 17153 3099 17187
rect 3893 17153 3927 17187
rect 2697 17085 2731 17119
rect 4077 17085 4111 17119
rect 3709 17017 3743 17051
rect 2973 16677 3007 16711
rect 1593 16609 1627 16643
rect 3065 16609 3099 16643
rect 5365 16609 5399 16643
rect 2789 16541 2823 16575
rect 2881 16541 2915 16575
rect 5098 16473 5132 16507
rect 3985 16405 4019 16439
rect 1685 16201 1719 16235
rect 5181 16201 5215 16235
rect 7941 16201 7975 16235
rect 4046 16133 4080 16167
rect 6806 16133 6840 16167
rect 1593 16065 1627 16099
rect 1869 16065 1903 16099
rect 2789 16065 2823 16099
rect 2973 16065 3007 16099
rect 3801 15997 3835 16031
rect 6561 15997 6595 16031
rect 2053 15861 2087 15895
rect 2789 15861 2823 15895
rect 1961 15657 1995 15691
rect 2789 15657 2823 15691
rect 7849 15657 7883 15691
rect 1593 15589 1627 15623
rect 2605 15589 2639 15623
rect 4629 15589 4663 15623
rect 6009 15453 6043 15487
rect 6469 15453 6503 15487
rect 1961 15385 1995 15419
rect 2757 15385 2791 15419
rect 2973 15385 3007 15419
rect 5742 15385 5776 15419
rect 6714 15385 6748 15419
rect 2145 15317 2179 15351
rect 2329 15113 2363 15147
rect 4261 15113 4295 15147
rect 7941 15113 7975 15147
rect 6828 15045 6862 15079
rect 3442 14977 3476 15011
rect 5549 14977 5583 15011
rect 3709 14909 3743 14943
rect 5825 14909 5859 14943
rect 6561 14909 6595 14943
rect 4169 14569 4203 14603
rect 5549 14365 5583 14399
rect 6193 14365 6227 14399
rect 6460 14365 6494 14399
rect 5282 14297 5316 14331
rect 7573 14229 7607 14263
rect 2690 14025 2724 14059
rect 5733 14025 5767 14059
rect 7941 14025 7975 14059
rect 2789 13957 2823 13991
rect 3341 13957 3375 13991
rect 2513 13889 2547 13923
rect 2605 13889 2639 13923
rect 3249 13889 3283 13923
rect 3433 13889 3467 13923
rect 4609 13889 4643 13923
rect 6828 13889 6862 13923
rect 4353 13821 4387 13855
rect 6561 13821 6595 13855
rect 2697 13481 2731 13515
rect 2973 13481 3007 13515
rect 2605 13345 2639 13379
rect 2789 13277 2823 13311
rect 2513 13209 2547 13243
rect 5273 13209 5307 13243
rect 6561 13141 6595 13175
rect 7941 12937 7975 12971
rect 6828 12869 6862 12903
rect 2145 12801 2179 12835
rect 4353 12801 4387 12835
rect 1869 12733 1903 12767
rect 6561 12733 6595 12767
rect 2053 12665 2087 12699
rect 1961 12597 1995 12631
rect 3065 12597 3099 12631
rect 7941 12393 7975 12427
rect 1593 12325 1627 12359
rect 5641 12257 5675 12291
rect 6561 12257 6595 12291
rect 1777 12189 1811 12223
rect 2421 12189 2455 12223
rect 2605 12189 2639 12223
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 3065 12121 3099 12155
rect 5374 12121 5408 12155
rect 6828 12121 6862 12155
rect 4261 12053 4295 12087
rect 2237 11849 2271 11883
rect 3065 11849 3099 11883
rect 1777 11781 1811 11815
rect 2145 11781 2179 11815
rect 2329 11713 2363 11747
rect 2973 11713 3007 11747
rect 3157 11713 3191 11747
rect 5098 11713 5132 11747
rect 5365 11713 5399 11747
rect 2513 11645 2547 11679
rect 3985 11577 4019 11611
rect 1777 11305 1811 11339
rect 7389 11305 7423 11339
rect 1593 11169 1627 11203
rect 6009 11169 6043 11203
rect 1869 11101 1903 11135
rect 1593 11033 1627 11067
rect 6254 11033 6288 11067
rect 7941 10761 7975 10795
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 5365 10217 5399 10251
rect 7113 10149 7147 10183
rect 3985 10081 4019 10115
rect 1593 10013 1627 10047
rect 4252 10013 4286 10047
rect 5825 9945 5859 9979
rect 1869 9605 1903 9639
rect 2069 9605 2103 9639
rect 6561 9605 6595 9639
rect 7941 9469 7975 9503
rect 8217 9469 8251 9503
rect 2053 9333 2087 9367
rect 2237 9333 2271 9367
rect 1961 8993 1995 9027
rect 1593 8925 1627 8959
rect 1685 8857 1719 8891
rect 1777 8789 1811 8823
rect 1961 8789 1995 8823
rect 2881 8585 2915 8619
rect 5181 8585 5215 8619
rect 2697 8517 2731 8551
rect 4068 8517 4102 8551
rect 2789 8449 2823 8483
rect 2329 8381 2363 8415
rect 3065 8381 3099 8415
rect 3801 8381 3835 8415
rect 2329 7905 2363 7939
rect 2145 7837 2179 7871
rect 1961 7701 1995 7735
rect 6653 7497 6687 7531
rect 7788 7429 7822 7463
rect 2237 7361 2271 7395
rect 2421 7361 2455 7395
rect 2513 7361 2547 7395
rect 8033 7361 8067 7395
rect 2329 7293 2363 7327
rect 2053 7157 2087 7191
rect 1685 6953 1719 6987
rect 2789 6817 2823 6851
rect 3985 6817 4019 6851
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 2421 6749 2455 6783
rect 2881 6749 2915 6783
rect 4252 6749 4286 6783
rect 1869 6681 1903 6715
rect 2513 6613 2547 6647
rect 2697 6613 2731 6647
rect 3065 6613 3099 6647
rect 5365 6613 5399 6647
rect 4629 6409 4663 6443
rect 7941 6409 7975 6443
rect 5764 6341 5798 6375
rect 2053 6273 2087 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2421 6273 2455 6307
rect 6009 6273 6043 6307
rect 6561 6273 6595 6307
rect 6828 6273 6862 6307
rect 2697 6069 2731 6103
rect 2513 5865 2547 5899
rect 6561 5865 6595 5899
rect 2605 5661 2639 5695
rect 5273 5661 5307 5695
rect 1593 5593 1627 5627
rect 1777 5593 1811 5627
rect 1961 5321 1995 5355
rect 3065 5321 3099 5355
rect 7941 5321 7975 5355
rect 4353 5253 4387 5287
rect 6828 5253 6862 5287
rect 1593 5185 1627 5219
rect 6561 5185 6595 5219
rect 2145 5049 2179 5083
rect 1961 4981 1995 5015
rect 2053 4777 2087 4811
rect 3433 4641 3467 4675
rect 4261 4641 4295 4675
rect 6193 4641 6227 4675
rect 3177 4573 3211 4607
rect 4528 4573 4562 4607
rect 6460 4573 6494 4607
rect 5641 4437 5675 4471
rect 7573 4437 7607 4471
rect 1961 4165 1995 4199
rect 1685 4097 1719 4131
rect 1777 4097 1811 4131
rect 2697 4097 2731 4131
rect 2881 4097 2915 4131
rect 5190 4097 5224 4131
rect 5457 4097 5491 4131
rect 6561 4097 6595 4131
rect 6837 4097 6871 4131
rect 2605 4029 2639 4063
rect 2789 4029 2823 4063
rect 7941 4029 7975 4063
rect 1961 3961 1995 3995
rect 4077 3961 4111 3995
rect 2421 3893 2455 3927
rect 2605 3689 2639 3723
rect 2789 3689 2823 3723
rect 7849 3689 7883 3723
rect 2237 3621 2271 3655
rect 3985 3553 4019 3587
rect 6285 3553 6319 3587
rect 6561 3553 6595 3587
rect 4252 3485 4286 3519
rect 2605 3417 2639 3451
rect 5365 3349 5399 3383
rect 2145 3145 2179 3179
rect 4252 3077 4286 3111
rect 1961 3009 1995 3043
rect 3985 3009 4019 3043
rect 1685 2941 1719 2975
rect 1777 2941 1811 2975
rect 1869 2941 1903 2975
rect 5365 2805 5399 2839
rect 1685 2601 1719 2635
rect 5365 2601 5399 2635
rect 2329 2465 2363 2499
rect 3985 2465 4019 2499
rect 15393 2465 15427 2499
rect 1593 2397 1627 2431
rect 1777 2397 1811 2431
rect 1869 2397 1903 2431
rect 4252 2397 4286 2431
rect 14933 2397 14967 2431
<< metal1 >>
rect 1104 47354 18860 47376
rect 1104 47302 3169 47354
rect 3221 47302 3233 47354
rect 3285 47302 3297 47354
rect 3349 47302 3361 47354
rect 3413 47302 3425 47354
rect 3477 47302 7608 47354
rect 7660 47302 7672 47354
rect 7724 47302 7736 47354
rect 7788 47302 7800 47354
rect 7852 47302 7864 47354
rect 7916 47302 12047 47354
rect 12099 47302 12111 47354
rect 12163 47302 12175 47354
rect 12227 47302 12239 47354
rect 12291 47302 12303 47354
rect 12355 47302 16486 47354
rect 16538 47302 16550 47354
rect 16602 47302 16614 47354
rect 16666 47302 16678 47354
rect 16730 47302 16742 47354
rect 16794 47302 18860 47354
rect 1104 47280 18860 47302
rect 934 47132 940 47184
rect 992 47172 998 47184
rect 1581 47175 1639 47181
rect 1581 47172 1593 47175
rect 992 47144 1593 47172
rect 992 47132 998 47144
rect 1581 47141 1593 47144
rect 1627 47141 1639 47175
rect 1581 47135 1639 47141
rect 1394 46928 1400 46980
rect 1452 46968 1458 46980
rect 1765 46971 1823 46977
rect 1765 46968 1777 46971
rect 1452 46940 1777 46968
rect 1452 46928 1458 46940
rect 1765 46937 1777 46940
rect 1811 46937 1823 46971
rect 1765 46931 1823 46937
rect 1104 46810 19019 46832
rect 1104 46758 5388 46810
rect 5440 46758 5452 46810
rect 5504 46758 5516 46810
rect 5568 46758 5580 46810
rect 5632 46758 5644 46810
rect 5696 46758 9827 46810
rect 9879 46758 9891 46810
rect 9943 46758 9955 46810
rect 10007 46758 10019 46810
rect 10071 46758 10083 46810
rect 10135 46758 14266 46810
rect 14318 46758 14330 46810
rect 14382 46758 14394 46810
rect 14446 46758 14458 46810
rect 14510 46758 14522 46810
rect 14574 46758 18705 46810
rect 18757 46758 18769 46810
rect 18821 46758 18833 46810
rect 18885 46758 18897 46810
rect 18949 46758 18961 46810
rect 19013 46758 19019 46810
rect 1104 46736 19019 46758
rect 1104 46266 18860 46288
rect 1104 46214 3169 46266
rect 3221 46214 3233 46266
rect 3285 46214 3297 46266
rect 3349 46214 3361 46266
rect 3413 46214 3425 46266
rect 3477 46214 7608 46266
rect 7660 46214 7672 46266
rect 7724 46214 7736 46266
rect 7788 46214 7800 46266
rect 7852 46214 7864 46266
rect 7916 46214 12047 46266
rect 12099 46214 12111 46266
rect 12163 46214 12175 46266
rect 12227 46214 12239 46266
rect 12291 46214 12303 46266
rect 12355 46214 16486 46266
rect 16538 46214 16550 46266
rect 16602 46214 16614 46266
rect 16666 46214 16678 46266
rect 16730 46214 16742 46266
rect 16794 46214 18860 46266
rect 1104 46192 18860 46214
rect 1104 45722 19019 45744
rect 1104 45670 5388 45722
rect 5440 45670 5452 45722
rect 5504 45670 5516 45722
rect 5568 45670 5580 45722
rect 5632 45670 5644 45722
rect 5696 45670 9827 45722
rect 9879 45670 9891 45722
rect 9943 45670 9955 45722
rect 10007 45670 10019 45722
rect 10071 45670 10083 45722
rect 10135 45670 14266 45722
rect 14318 45670 14330 45722
rect 14382 45670 14394 45722
rect 14446 45670 14458 45722
rect 14510 45670 14522 45722
rect 14574 45670 18705 45722
rect 18757 45670 18769 45722
rect 18821 45670 18833 45722
rect 18885 45670 18897 45722
rect 18949 45670 18961 45722
rect 19013 45670 19019 45722
rect 1104 45648 19019 45670
rect 1104 45178 18860 45200
rect 1104 45126 3169 45178
rect 3221 45126 3233 45178
rect 3285 45126 3297 45178
rect 3349 45126 3361 45178
rect 3413 45126 3425 45178
rect 3477 45126 7608 45178
rect 7660 45126 7672 45178
rect 7724 45126 7736 45178
rect 7788 45126 7800 45178
rect 7852 45126 7864 45178
rect 7916 45126 12047 45178
rect 12099 45126 12111 45178
rect 12163 45126 12175 45178
rect 12227 45126 12239 45178
rect 12291 45126 12303 45178
rect 12355 45126 16486 45178
rect 16538 45126 16550 45178
rect 16602 45126 16614 45178
rect 16666 45126 16678 45178
rect 16730 45126 16742 45178
rect 16794 45126 18860 45178
rect 1104 45104 18860 45126
rect 934 44820 940 44872
rect 992 44860 998 44872
rect 1581 44863 1639 44869
rect 1581 44860 1593 44863
rect 992 44832 1593 44860
rect 992 44820 998 44832
rect 1581 44829 1593 44832
rect 1627 44829 1639 44863
rect 1581 44823 1639 44829
rect 1104 44634 19019 44656
rect 1104 44582 5388 44634
rect 5440 44582 5452 44634
rect 5504 44582 5516 44634
rect 5568 44582 5580 44634
rect 5632 44582 5644 44634
rect 5696 44582 9827 44634
rect 9879 44582 9891 44634
rect 9943 44582 9955 44634
rect 10007 44582 10019 44634
rect 10071 44582 10083 44634
rect 10135 44582 14266 44634
rect 14318 44582 14330 44634
rect 14382 44582 14394 44634
rect 14446 44582 14458 44634
rect 14510 44582 14522 44634
rect 14574 44582 18705 44634
rect 18757 44582 18769 44634
rect 18821 44582 18833 44634
rect 18885 44582 18897 44634
rect 18949 44582 18961 44634
rect 19013 44582 19019 44634
rect 1104 44560 19019 44582
rect 1104 44090 18860 44112
rect 1104 44038 3169 44090
rect 3221 44038 3233 44090
rect 3285 44038 3297 44090
rect 3349 44038 3361 44090
rect 3413 44038 3425 44090
rect 3477 44038 7608 44090
rect 7660 44038 7672 44090
rect 7724 44038 7736 44090
rect 7788 44038 7800 44090
rect 7852 44038 7864 44090
rect 7916 44038 12047 44090
rect 12099 44038 12111 44090
rect 12163 44038 12175 44090
rect 12227 44038 12239 44090
rect 12291 44038 12303 44090
rect 12355 44038 16486 44090
rect 16538 44038 16550 44090
rect 16602 44038 16614 44090
rect 16666 44038 16678 44090
rect 16730 44038 16742 44090
rect 16794 44038 18860 44090
rect 1104 44016 18860 44038
rect 1104 43546 19019 43568
rect 1104 43494 5388 43546
rect 5440 43494 5452 43546
rect 5504 43494 5516 43546
rect 5568 43494 5580 43546
rect 5632 43494 5644 43546
rect 5696 43494 9827 43546
rect 9879 43494 9891 43546
rect 9943 43494 9955 43546
rect 10007 43494 10019 43546
rect 10071 43494 10083 43546
rect 10135 43494 14266 43546
rect 14318 43494 14330 43546
rect 14382 43494 14394 43546
rect 14446 43494 14458 43546
rect 14510 43494 14522 43546
rect 14574 43494 18705 43546
rect 18757 43494 18769 43546
rect 18821 43494 18833 43546
rect 18885 43494 18897 43546
rect 18949 43494 18961 43546
rect 19013 43494 19019 43546
rect 1104 43472 19019 43494
rect 1104 43002 18860 43024
rect 1104 42950 3169 43002
rect 3221 42950 3233 43002
rect 3285 42950 3297 43002
rect 3349 42950 3361 43002
rect 3413 42950 3425 43002
rect 3477 42950 7608 43002
rect 7660 42950 7672 43002
rect 7724 42950 7736 43002
rect 7788 42950 7800 43002
rect 7852 42950 7864 43002
rect 7916 42950 12047 43002
rect 12099 42950 12111 43002
rect 12163 42950 12175 43002
rect 12227 42950 12239 43002
rect 12291 42950 12303 43002
rect 12355 42950 16486 43002
rect 16538 42950 16550 43002
rect 16602 42950 16614 43002
rect 16666 42950 16678 43002
rect 16730 42950 16742 43002
rect 16794 42950 18860 43002
rect 1104 42928 18860 42950
rect 1104 42458 19019 42480
rect 1104 42406 5388 42458
rect 5440 42406 5452 42458
rect 5504 42406 5516 42458
rect 5568 42406 5580 42458
rect 5632 42406 5644 42458
rect 5696 42406 9827 42458
rect 9879 42406 9891 42458
rect 9943 42406 9955 42458
rect 10007 42406 10019 42458
rect 10071 42406 10083 42458
rect 10135 42406 14266 42458
rect 14318 42406 14330 42458
rect 14382 42406 14394 42458
rect 14446 42406 14458 42458
rect 14510 42406 14522 42458
rect 14574 42406 18705 42458
rect 18757 42406 18769 42458
rect 18821 42406 18833 42458
rect 18885 42406 18897 42458
rect 18949 42406 18961 42458
rect 19013 42406 19019 42458
rect 1104 42384 19019 42406
rect 1104 41914 18860 41936
rect 1104 41862 3169 41914
rect 3221 41862 3233 41914
rect 3285 41862 3297 41914
rect 3349 41862 3361 41914
rect 3413 41862 3425 41914
rect 3477 41862 7608 41914
rect 7660 41862 7672 41914
rect 7724 41862 7736 41914
rect 7788 41862 7800 41914
rect 7852 41862 7864 41914
rect 7916 41862 12047 41914
rect 12099 41862 12111 41914
rect 12163 41862 12175 41914
rect 12227 41862 12239 41914
rect 12291 41862 12303 41914
rect 12355 41862 16486 41914
rect 16538 41862 16550 41914
rect 16602 41862 16614 41914
rect 16666 41862 16678 41914
rect 16730 41862 16742 41914
rect 16794 41862 18860 41914
rect 1104 41840 18860 41862
rect 1104 41370 19019 41392
rect 1104 41318 5388 41370
rect 5440 41318 5452 41370
rect 5504 41318 5516 41370
rect 5568 41318 5580 41370
rect 5632 41318 5644 41370
rect 5696 41318 9827 41370
rect 9879 41318 9891 41370
rect 9943 41318 9955 41370
rect 10007 41318 10019 41370
rect 10071 41318 10083 41370
rect 10135 41318 14266 41370
rect 14318 41318 14330 41370
rect 14382 41318 14394 41370
rect 14446 41318 14458 41370
rect 14510 41318 14522 41370
rect 14574 41318 18705 41370
rect 18757 41318 18769 41370
rect 18821 41318 18833 41370
rect 18885 41318 18897 41370
rect 18949 41318 18961 41370
rect 19013 41318 19019 41370
rect 1104 41296 19019 41318
rect 1765 41123 1823 41129
rect 1765 41089 1777 41123
rect 1811 41120 1823 41123
rect 2498 41120 2504 41132
rect 1811 41092 2504 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 2498 41080 2504 41092
rect 2556 41080 2562 41132
rect 934 40944 940 40996
rect 992 40984 998 40996
rect 1581 40987 1639 40993
rect 1581 40984 1593 40987
rect 992 40956 1593 40984
rect 992 40944 998 40956
rect 1581 40953 1593 40956
rect 1627 40953 1639 40987
rect 1581 40947 1639 40953
rect 1104 40826 18860 40848
rect 1104 40774 3169 40826
rect 3221 40774 3233 40826
rect 3285 40774 3297 40826
rect 3349 40774 3361 40826
rect 3413 40774 3425 40826
rect 3477 40774 7608 40826
rect 7660 40774 7672 40826
rect 7724 40774 7736 40826
rect 7788 40774 7800 40826
rect 7852 40774 7864 40826
rect 7916 40774 12047 40826
rect 12099 40774 12111 40826
rect 12163 40774 12175 40826
rect 12227 40774 12239 40826
rect 12291 40774 12303 40826
rect 12355 40774 16486 40826
rect 16538 40774 16550 40826
rect 16602 40774 16614 40826
rect 16666 40774 16678 40826
rect 16730 40774 16742 40826
rect 16794 40774 18860 40826
rect 1104 40752 18860 40774
rect 1104 40282 19019 40304
rect 1104 40230 5388 40282
rect 5440 40230 5452 40282
rect 5504 40230 5516 40282
rect 5568 40230 5580 40282
rect 5632 40230 5644 40282
rect 5696 40230 9827 40282
rect 9879 40230 9891 40282
rect 9943 40230 9955 40282
rect 10007 40230 10019 40282
rect 10071 40230 10083 40282
rect 10135 40230 14266 40282
rect 14318 40230 14330 40282
rect 14382 40230 14394 40282
rect 14446 40230 14458 40282
rect 14510 40230 14522 40282
rect 14574 40230 18705 40282
rect 18757 40230 18769 40282
rect 18821 40230 18833 40282
rect 18885 40230 18897 40282
rect 18949 40230 18961 40282
rect 19013 40230 19019 40282
rect 1104 40208 19019 40230
rect 1104 39738 18860 39760
rect 1104 39686 3169 39738
rect 3221 39686 3233 39738
rect 3285 39686 3297 39738
rect 3349 39686 3361 39738
rect 3413 39686 3425 39738
rect 3477 39686 7608 39738
rect 7660 39686 7672 39738
rect 7724 39686 7736 39738
rect 7788 39686 7800 39738
rect 7852 39686 7864 39738
rect 7916 39686 12047 39738
rect 12099 39686 12111 39738
rect 12163 39686 12175 39738
rect 12227 39686 12239 39738
rect 12291 39686 12303 39738
rect 12355 39686 16486 39738
rect 16538 39686 16550 39738
rect 16602 39686 16614 39738
rect 16666 39686 16678 39738
rect 16730 39686 16742 39738
rect 16794 39686 18860 39738
rect 1104 39664 18860 39686
rect 1104 39194 19019 39216
rect 1104 39142 5388 39194
rect 5440 39142 5452 39194
rect 5504 39142 5516 39194
rect 5568 39142 5580 39194
rect 5632 39142 5644 39194
rect 5696 39142 9827 39194
rect 9879 39142 9891 39194
rect 9943 39142 9955 39194
rect 10007 39142 10019 39194
rect 10071 39142 10083 39194
rect 10135 39142 14266 39194
rect 14318 39142 14330 39194
rect 14382 39142 14394 39194
rect 14446 39142 14458 39194
rect 14510 39142 14522 39194
rect 14574 39142 18705 39194
rect 18757 39142 18769 39194
rect 18821 39142 18833 39194
rect 18885 39142 18897 39194
rect 18949 39142 18961 39194
rect 19013 39142 19019 39194
rect 1104 39120 19019 39142
rect 1104 38650 18860 38672
rect 1104 38598 3169 38650
rect 3221 38598 3233 38650
rect 3285 38598 3297 38650
rect 3349 38598 3361 38650
rect 3413 38598 3425 38650
rect 3477 38598 7608 38650
rect 7660 38598 7672 38650
rect 7724 38598 7736 38650
rect 7788 38598 7800 38650
rect 7852 38598 7864 38650
rect 7916 38598 12047 38650
rect 12099 38598 12111 38650
rect 12163 38598 12175 38650
rect 12227 38598 12239 38650
rect 12291 38598 12303 38650
rect 12355 38598 16486 38650
rect 16538 38598 16550 38650
rect 16602 38598 16614 38650
rect 16666 38598 16678 38650
rect 16730 38598 16742 38650
rect 16794 38598 18860 38650
rect 1104 38576 18860 38598
rect 1104 38106 19019 38128
rect 1104 38054 5388 38106
rect 5440 38054 5452 38106
rect 5504 38054 5516 38106
rect 5568 38054 5580 38106
rect 5632 38054 5644 38106
rect 5696 38054 9827 38106
rect 9879 38054 9891 38106
rect 9943 38054 9955 38106
rect 10007 38054 10019 38106
rect 10071 38054 10083 38106
rect 10135 38054 14266 38106
rect 14318 38054 14330 38106
rect 14382 38054 14394 38106
rect 14446 38054 14458 38106
rect 14510 38054 14522 38106
rect 14574 38054 18705 38106
rect 18757 38054 18769 38106
rect 18821 38054 18833 38106
rect 18885 38054 18897 38106
rect 18949 38054 18961 38106
rect 19013 38054 19019 38106
rect 1104 38032 19019 38054
rect 934 37612 940 37664
rect 992 37652 998 37664
rect 1581 37655 1639 37661
rect 1581 37652 1593 37655
rect 992 37624 1593 37652
rect 992 37612 998 37624
rect 1581 37621 1593 37624
rect 1627 37621 1639 37655
rect 1581 37615 1639 37621
rect 1104 37562 18860 37584
rect 1104 37510 3169 37562
rect 3221 37510 3233 37562
rect 3285 37510 3297 37562
rect 3349 37510 3361 37562
rect 3413 37510 3425 37562
rect 3477 37510 7608 37562
rect 7660 37510 7672 37562
rect 7724 37510 7736 37562
rect 7788 37510 7800 37562
rect 7852 37510 7864 37562
rect 7916 37510 12047 37562
rect 12099 37510 12111 37562
rect 12163 37510 12175 37562
rect 12227 37510 12239 37562
rect 12291 37510 12303 37562
rect 12355 37510 16486 37562
rect 16538 37510 16550 37562
rect 16602 37510 16614 37562
rect 16666 37510 16678 37562
rect 16730 37510 16742 37562
rect 16794 37510 18860 37562
rect 1104 37488 18860 37510
rect 1104 37018 19019 37040
rect 1104 36966 5388 37018
rect 5440 36966 5452 37018
rect 5504 36966 5516 37018
rect 5568 36966 5580 37018
rect 5632 36966 5644 37018
rect 5696 36966 9827 37018
rect 9879 36966 9891 37018
rect 9943 36966 9955 37018
rect 10007 36966 10019 37018
rect 10071 36966 10083 37018
rect 10135 36966 14266 37018
rect 14318 36966 14330 37018
rect 14382 36966 14394 37018
rect 14446 36966 14458 37018
rect 14510 36966 14522 37018
rect 14574 36966 18705 37018
rect 18757 36966 18769 37018
rect 18821 36966 18833 37018
rect 18885 36966 18897 37018
rect 18949 36966 18961 37018
rect 19013 36966 19019 37018
rect 1104 36944 19019 36966
rect 1104 36474 18860 36496
rect 1104 36422 3169 36474
rect 3221 36422 3233 36474
rect 3285 36422 3297 36474
rect 3349 36422 3361 36474
rect 3413 36422 3425 36474
rect 3477 36422 7608 36474
rect 7660 36422 7672 36474
rect 7724 36422 7736 36474
rect 7788 36422 7800 36474
rect 7852 36422 7864 36474
rect 7916 36422 12047 36474
rect 12099 36422 12111 36474
rect 12163 36422 12175 36474
rect 12227 36422 12239 36474
rect 12291 36422 12303 36474
rect 12355 36422 16486 36474
rect 16538 36422 16550 36474
rect 16602 36422 16614 36474
rect 16666 36422 16678 36474
rect 16730 36422 16742 36474
rect 16794 36422 18860 36474
rect 1104 36400 18860 36422
rect 6825 36227 6883 36233
rect 6825 36193 6837 36227
rect 6871 36224 6883 36227
rect 7282 36224 7288 36236
rect 6871 36196 7288 36224
rect 6871 36193 6883 36196
rect 6825 36187 6883 36193
rect 7282 36184 7288 36196
rect 7340 36184 7346 36236
rect 6365 36159 6423 36165
rect 6365 36125 6377 36159
rect 6411 36125 6423 36159
rect 6365 36119 6423 36125
rect 6733 36159 6791 36165
rect 6733 36125 6745 36159
rect 6779 36156 6791 36159
rect 7190 36156 7196 36168
rect 6779 36128 7196 36156
rect 6779 36125 6791 36128
rect 6733 36119 6791 36125
rect 4614 36048 4620 36100
rect 4672 36088 4678 36100
rect 5905 36091 5963 36097
rect 5905 36088 5917 36091
rect 4672 36060 5917 36088
rect 4672 36048 4678 36060
rect 5905 36057 5917 36060
rect 5951 36057 5963 36091
rect 6380 36088 6408 36119
rect 7190 36116 7196 36128
rect 7248 36116 7254 36168
rect 6914 36088 6920 36100
rect 6380 36060 6920 36088
rect 5905 36051 5963 36057
rect 6914 36048 6920 36060
rect 6972 36048 6978 36100
rect 1104 35930 19019 35952
rect 1104 35878 5388 35930
rect 5440 35878 5452 35930
rect 5504 35878 5516 35930
rect 5568 35878 5580 35930
rect 5632 35878 5644 35930
rect 5696 35878 9827 35930
rect 9879 35878 9891 35930
rect 9943 35878 9955 35930
rect 10007 35878 10019 35930
rect 10071 35878 10083 35930
rect 10135 35878 14266 35930
rect 14318 35878 14330 35930
rect 14382 35878 14394 35930
rect 14446 35878 14458 35930
rect 14510 35878 14522 35930
rect 14574 35878 18705 35930
rect 18757 35878 18769 35930
rect 18821 35878 18833 35930
rect 18885 35878 18897 35930
rect 18949 35878 18961 35930
rect 19013 35878 19019 35930
rect 1104 35856 19019 35878
rect 4614 35640 4620 35692
rect 4672 35640 4678 35692
rect 4801 35683 4859 35689
rect 4801 35649 4813 35683
rect 4847 35680 4859 35683
rect 6178 35680 6184 35692
rect 4847 35652 6184 35680
rect 4847 35649 4859 35652
rect 4801 35643 4859 35649
rect 6178 35640 6184 35652
rect 6236 35640 6242 35692
rect 4709 35479 4767 35485
rect 4709 35445 4721 35479
rect 4755 35476 4767 35479
rect 5258 35476 5264 35488
rect 4755 35448 5264 35476
rect 4755 35445 4767 35448
rect 4709 35439 4767 35445
rect 5258 35436 5264 35448
rect 5316 35436 5322 35488
rect 1104 35386 18860 35408
rect 1104 35334 3169 35386
rect 3221 35334 3233 35386
rect 3285 35334 3297 35386
rect 3349 35334 3361 35386
rect 3413 35334 3425 35386
rect 3477 35334 7608 35386
rect 7660 35334 7672 35386
rect 7724 35334 7736 35386
rect 7788 35334 7800 35386
rect 7852 35334 7864 35386
rect 7916 35334 12047 35386
rect 12099 35334 12111 35386
rect 12163 35334 12175 35386
rect 12227 35334 12239 35386
rect 12291 35334 12303 35386
rect 12355 35334 16486 35386
rect 16538 35334 16550 35386
rect 16602 35334 16614 35386
rect 16666 35334 16678 35386
rect 16730 35334 16742 35386
rect 16794 35334 18860 35386
rect 1104 35312 18860 35334
rect 6086 35028 6092 35080
rect 6144 35028 6150 35080
rect 6914 35028 6920 35080
rect 6972 35028 6978 35080
rect 6362 34892 6368 34944
rect 6420 34892 6426 34944
rect 1104 34842 19019 34864
rect 1104 34790 5388 34842
rect 5440 34790 5452 34842
rect 5504 34790 5516 34842
rect 5568 34790 5580 34842
rect 5632 34790 5644 34842
rect 5696 34790 9827 34842
rect 9879 34790 9891 34842
rect 9943 34790 9955 34842
rect 10007 34790 10019 34842
rect 10071 34790 10083 34842
rect 10135 34790 14266 34842
rect 14318 34790 14330 34842
rect 14382 34790 14394 34842
rect 14446 34790 14458 34842
rect 14510 34790 14522 34842
rect 14574 34790 18705 34842
rect 18757 34790 18769 34842
rect 18821 34790 18833 34842
rect 18885 34790 18897 34842
rect 18949 34790 18961 34842
rect 19013 34790 19019 34842
rect 1104 34768 19019 34790
rect 6914 34620 6920 34672
rect 6972 34660 6978 34672
rect 6972 34632 7512 34660
rect 6972 34620 6978 34632
rect 6454 34552 6460 34604
rect 6512 34592 6518 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 6512 34564 6561 34592
rect 6512 34552 6518 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 6549 34555 6607 34561
rect 7282 34552 7288 34604
rect 7340 34552 7346 34604
rect 7484 34601 7512 34632
rect 7469 34595 7527 34601
rect 7469 34561 7481 34595
rect 7515 34561 7527 34595
rect 7469 34555 7527 34561
rect 6178 34348 6184 34400
rect 6236 34388 6242 34400
rect 6733 34391 6791 34397
rect 6733 34388 6745 34391
rect 6236 34360 6745 34388
rect 6236 34348 6242 34360
rect 6733 34357 6745 34360
rect 6779 34357 6791 34391
rect 6733 34351 6791 34357
rect 1104 34298 18860 34320
rect 1104 34246 3169 34298
rect 3221 34246 3233 34298
rect 3285 34246 3297 34298
rect 3349 34246 3361 34298
rect 3413 34246 3425 34298
rect 3477 34246 7608 34298
rect 7660 34246 7672 34298
rect 7724 34246 7736 34298
rect 7788 34246 7800 34298
rect 7852 34246 7864 34298
rect 7916 34246 12047 34298
rect 12099 34246 12111 34298
rect 12163 34246 12175 34298
rect 12227 34246 12239 34298
rect 12291 34246 12303 34298
rect 12355 34246 16486 34298
rect 16538 34246 16550 34298
rect 16602 34246 16614 34298
rect 16666 34246 16678 34298
rect 16730 34246 16742 34298
rect 16794 34246 18860 34298
rect 1104 34224 18860 34246
rect 6273 34187 6331 34193
rect 6273 34153 6285 34187
rect 6319 34184 6331 34187
rect 6362 34184 6368 34196
rect 6319 34156 6368 34184
rect 6319 34153 6331 34156
rect 6273 34147 6331 34153
rect 6362 34144 6368 34156
rect 6420 34144 6426 34196
rect 7374 34144 7380 34196
rect 7432 34184 7438 34196
rect 7561 34187 7619 34193
rect 7561 34184 7573 34187
rect 7432 34156 7573 34184
rect 7432 34144 7438 34156
rect 7561 34153 7573 34156
rect 7607 34153 7619 34187
rect 7561 34147 7619 34153
rect 6825 34119 6883 34125
rect 6825 34085 6837 34119
rect 6871 34116 6883 34119
rect 8662 34116 8668 34128
rect 6871 34088 8668 34116
rect 6871 34085 6883 34088
rect 6825 34079 6883 34085
rect 8662 34076 8668 34088
rect 8720 34076 8726 34128
rect 5718 34008 5724 34060
rect 5776 34048 5782 34060
rect 6178 34048 6184 34060
rect 5776 34020 6184 34048
rect 5776 34008 5782 34020
rect 6178 34008 6184 34020
rect 6236 34008 6242 34060
rect 7190 34008 7196 34060
rect 7248 34048 7254 34060
rect 7248 34020 7696 34048
rect 7248 34008 7254 34020
rect 6454 33940 6460 33992
rect 6512 33980 6518 33992
rect 6643 33983 6701 33989
rect 6643 33980 6655 33983
rect 6512 33952 6655 33980
rect 6512 33940 6518 33952
rect 6643 33949 6655 33952
rect 6689 33949 6701 33983
rect 6643 33943 6701 33949
rect 7282 33940 7288 33992
rect 7340 33980 7346 33992
rect 7340 33952 7604 33980
rect 7340 33940 7346 33952
rect 934 33872 940 33924
rect 992 33912 998 33924
rect 1581 33915 1639 33921
rect 1581 33912 1593 33915
rect 992 33884 1593 33912
rect 992 33872 998 33884
rect 1581 33881 1593 33884
rect 1627 33881 1639 33915
rect 1581 33875 1639 33881
rect 1670 33872 1676 33924
rect 1728 33912 1734 33924
rect 7576 33921 7604 33952
rect 1765 33915 1823 33921
rect 1765 33912 1777 33915
rect 1728 33884 1777 33912
rect 1728 33872 1734 33884
rect 1765 33881 1777 33884
rect 1811 33881 1823 33915
rect 1765 33875 1823 33881
rect 7545 33915 7604 33921
rect 7545 33881 7557 33915
rect 7591 33884 7604 33915
rect 7668 33912 7696 34020
rect 7745 33915 7803 33921
rect 7745 33912 7757 33915
rect 7668 33884 7757 33912
rect 7591 33881 7603 33884
rect 7545 33875 7603 33881
rect 7745 33881 7757 33884
rect 7791 33881 7803 33915
rect 7745 33875 7803 33881
rect 6641 33847 6699 33853
rect 6641 33813 6653 33847
rect 6687 33844 6699 33847
rect 7377 33847 7435 33853
rect 7377 33844 7389 33847
rect 6687 33816 7389 33844
rect 6687 33813 6699 33816
rect 6641 33807 6699 33813
rect 7377 33813 7389 33816
rect 7423 33813 7435 33847
rect 7377 33807 7435 33813
rect 1104 33754 19019 33776
rect 1104 33702 5388 33754
rect 5440 33702 5452 33754
rect 5504 33702 5516 33754
rect 5568 33702 5580 33754
rect 5632 33702 5644 33754
rect 5696 33702 9827 33754
rect 9879 33702 9891 33754
rect 9943 33702 9955 33754
rect 10007 33702 10019 33754
rect 10071 33702 10083 33754
rect 10135 33702 14266 33754
rect 14318 33702 14330 33754
rect 14382 33702 14394 33754
rect 14446 33702 14458 33754
rect 14510 33702 14522 33754
rect 14574 33702 18705 33754
rect 18757 33702 18769 33754
rect 18821 33702 18833 33754
rect 18885 33702 18897 33754
rect 18949 33702 18961 33754
rect 19013 33702 19019 33754
rect 1104 33680 19019 33702
rect 1104 33210 18860 33232
rect 1104 33158 3169 33210
rect 3221 33158 3233 33210
rect 3285 33158 3297 33210
rect 3349 33158 3361 33210
rect 3413 33158 3425 33210
rect 3477 33158 7608 33210
rect 7660 33158 7672 33210
rect 7724 33158 7736 33210
rect 7788 33158 7800 33210
rect 7852 33158 7864 33210
rect 7916 33158 12047 33210
rect 12099 33158 12111 33210
rect 12163 33158 12175 33210
rect 12227 33158 12239 33210
rect 12291 33158 12303 33210
rect 12355 33158 16486 33210
rect 16538 33158 16550 33210
rect 16602 33158 16614 33210
rect 16666 33158 16678 33210
rect 16730 33158 16742 33210
rect 16794 33158 18860 33210
rect 1104 33136 18860 33158
rect 7190 33056 7196 33108
rect 7248 33096 7254 33108
rect 7285 33099 7343 33105
rect 7285 33096 7297 33099
rect 7248 33068 7297 33096
rect 7248 33056 7254 33068
rect 7285 33065 7297 33068
rect 7331 33065 7343 33099
rect 7285 33059 7343 33065
rect 5445 33031 5503 33037
rect 5445 32997 5457 33031
rect 5491 33028 5503 33031
rect 6086 33028 6092 33040
rect 5491 33000 6092 33028
rect 5491 32997 5503 33000
rect 5445 32991 5503 32997
rect 6086 32988 6092 33000
rect 6144 32988 6150 33040
rect 6178 32988 6184 33040
rect 6236 33028 6242 33040
rect 6236 33000 6914 33028
rect 6236 32988 6242 33000
rect 6886 32960 6914 33000
rect 7469 32963 7527 32969
rect 7469 32960 7481 32963
rect 6886 32932 7481 32960
rect 7469 32929 7481 32932
rect 7515 32929 7527 32963
rect 7469 32923 7527 32929
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32892 5779 32895
rect 6178 32892 6184 32904
rect 5767 32864 6184 32892
rect 5767 32861 5779 32864
rect 5721 32855 5779 32861
rect 6178 32852 6184 32864
rect 6236 32852 6242 32904
rect 6365 32895 6423 32901
rect 6365 32861 6377 32895
rect 6411 32861 6423 32895
rect 7098 32892 7104 32904
rect 6365 32855 6423 32861
rect 6886 32864 7104 32892
rect 6380 32824 6408 32855
rect 6886 32824 6914 32864
rect 7098 32852 7104 32864
rect 7156 32892 7162 32904
rect 7561 32895 7619 32901
rect 7561 32892 7573 32895
rect 7156 32864 7573 32892
rect 7156 32852 7162 32864
rect 7561 32861 7573 32864
rect 7607 32861 7619 32895
rect 7561 32855 7619 32861
rect 6380 32796 6914 32824
rect 7926 32716 7932 32768
rect 7984 32716 7990 32768
rect 1104 32666 19019 32688
rect 1104 32614 5388 32666
rect 5440 32614 5452 32666
rect 5504 32614 5516 32666
rect 5568 32614 5580 32666
rect 5632 32614 5644 32666
rect 5696 32614 9827 32666
rect 9879 32614 9891 32666
rect 9943 32614 9955 32666
rect 10007 32614 10019 32666
rect 10071 32614 10083 32666
rect 10135 32614 14266 32666
rect 14318 32614 14330 32666
rect 14382 32614 14394 32666
rect 14446 32614 14458 32666
rect 14510 32614 14522 32666
rect 14574 32614 18705 32666
rect 18757 32614 18769 32666
rect 18821 32614 18833 32666
rect 18885 32614 18897 32666
rect 18949 32614 18961 32666
rect 19013 32614 19019 32666
rect 1104 32592 19019 32614
rect 5718 32484 5724 32496
rect 5368 32456 5724 32484
rect 4614 32376 4620 32428
rect 4672 32416 4678 32428
rect 5166 32416 5172 32428
rect 4672 32388 5172 32416
rect 4672 32376 4678 32388
rect 5166 32376 5172 32388
rect 5224 32376 5230 32428
rect 5368 32425 5396 32456
rect 5718 32444 5724 32456
rect 5776 32444 5782 32496
rect 5353 32419 5411 32425
rect 5353 32385 5365 32419
rect 5399 32385 5411 32419
rect 5353 32379 5411 32385
rect 5445 32419 5503 32425
rect 5445 32385 5457 32419
rect 5491 32385 5503 32419
rect 5445 32379 5503 32385
rect 5537 32419 5595 32425
rect 5537 32385 5549 32419
rect 5583 32416 5595 32419
rect 6822 32416 6828 32428
rect 5583 32388 6828 32416
rect 5583 32385 5595 32388
rect 5537 32379 5595 32385
rect 5460 32280 5488 32379
rect 6822 32376 6828 32388
rect 6880 32416 6886 32428
rect 6914 32416 6920 32428
rect 6880 32388 6920 32416
rect 6880 32376 6886 32388
rect 6914 32376 6920 32388
rect 6972 32376 6978 32428
rect 6086 32280 6092 32292
rect 5460 32252 6092 32280
rect 6086 32240 6092 32252
rect 6144 32240 6150 32292
rect 5813 32215 5871 32221
rect 5813 32181 5825 32215
rect 5859 32212 5871 32215
rect 6638 32212 6644 32224
rect 5859 32184 6644 32212
rect 5859 32181 5871 32184
rect 5813 32175 5871 32181
rect 6638 32172 6644 32184
rect 6696 32172 6702 32224
rect 1104 32122 18860 32144
rect 1104 32070 3169 32122
rect 3221 32070 3233 32122
rect 3285 32070 3297 32122
rect 3349 32070 3361 32122
rect 3413 32070 3425 32122
rect 3477 32070 7608 32122
rect 7660 32070 7672 32122
rect 7724 32070 7736 32122
rect 7788 32070 7800 32122
rect 7852 32070 7864 32122
rect 7916 32070 12047 32122
rect 12099 32070 12111 32122
rect 12163 32070 12175 32122
rect 12227 32070 12239 32122
rect 12291 32070 12303 32122
rect 12355 32070 16486 32122
rect 16538 32070 16550 32122
rect 16602 32070 16614 32122
rect 16666 32070 16678 32122
rect 16730 32070 16742 32122
rect 16794 32070 18860 32122
rect 1104 32048 18860 32070
rect 5258 31764 5264 31816
rect 5316 31764 5322 31816
rect 5902 31764 5908 31816
rect 5960 31764 5966 31816
rect 4706 31696 4712 31748
rect 4764 31696 4770 31748
rect 1104 31578 19019 31600
rect 1104 31526 5388 31578
rect 5440 31526 5452 31578
rect 5504 31526 5516 31578
rect 5568 31526 5580 31578
rect 5632 31526 5644 31578
rect 5696 31526 9827 31578
rect 9879 31526 9891 31578
rect 9943 31526 9955 31578
rect 10007 31526 10019 31578
rect 10071 31526 10083 31578
rect 10135 31526 14266 31578
rect 14318 31526 14330 31578
rect 14382 31526 14394 31578
rect 14446 31526 14458 31578
rect 14510 31526 14522 31578
rect 14574 31526 18705 31578
rect 18757 31526 18769 31578
rect 18821 31526 18833 31578
rect 18885 31526 18897 31578
rect 18949 31526 18961 31578
rect 19013 31526 19019 31578
rect 1104 31504 19019 31526
rect 5902 31424 5908 31476
rect 5960 31464 5966 31476
rect 5960 31436 6776 31464
rect 5960 31424 5966 31436
rect 6454 31396 6460 31408
rect 5644 31368 6460 31396
rect 5644 31340 5672 31368
rect 6454 31356 6460 31368
rect 6512 31356 6518 31408
rect 5445 31331 5503 31337
rect 5445 31297 5457 31331
rect 5491 31328 5503 31331
rect 5626 31328 5632 31340
rect 5491 31300 5632 31328
rect 5491 31297 5503 31300
rect 5445 31291 5503 31297
rect 5626 31288 5632 31300
rect 5684 31288 5690 31340
rect 5994 31288 6000 31340
rect 6052 31328 6058 31340
rect 6362 31328 6368 31340
rect 6052 31300 6368 31328
rect 6052 31288 6058 31300
rect 6362 31288 6368 31300
rect 6420 31288 6426 31340
rect 6748 31337 6776 31436
rect 6733 31331 6791 31337
rect 6733 31297 6745 31331
rect 6779 31297 6791 31331
rect 6733 31291 6791 31297
rect 6822 31288 6828 31340
rect 6880 31288 6886 31340
rect 7009 31331 7067 31337
rect 7009 31297 7021 31331
rect 7055 31297 7067 31331
rect 7009 31291 7067 31297
rect 5166 31220 5172 31272
rect 5224 31260 5230 31272
rect 6840 31260 6868 31288
rect 5224 31232 6868 31260
rect 7024 31260 7052 31291
rect 7098 31288 7104 31340
rect 7156 31288 7162 31340
rect 7282 31260 7288 31272
rect 7024 31232 7288 31260
rect 5224 31220 5230 31232
rect 7282 31220 7288 31232
rect 7340 31220 7346 31272
rect 6549 31127 6607 31133
rect 6549 31093 6561 31127
rect 6595 31124 6607 31127
rect 8846 31124 8852 31136
rect 6595 31096 8852 31124
rect 6595 31093 6607 31096
rect 6549 31087 6607 31093
rect 8846 31084 8852 31096
rect 8904 31084 8910 31136
rect 1104 31034 18860 31056
rect 1104 30982 3169 31034
rect 3221 30982 3233 31034
rect 3285 30982 3297 31034
rect 3349 30982 3361 31034
rect 3413 30982 3425 31034
rect 3477 30982 7608 31034
rect 7660 30982 7672 31034
rect 7724 30982 7736 31034
rect 7788 30982 7800 31034
rect 7852 30982 7864 31034
rect 7916 30982 12047 31034
rect 12099 30982 12111 31034
rect 12163 30982 12175 31034
rect 12227 30982 12239 31034
rect 12291 30982 12303 31034
rect 12355 30982 16486 31034
rect 16538 30982 16550 31034
rect 16602 30982 16614 31034
rect 16666 30982 16678 31034
rect 16730 30982 16742 31034
rect 16794 30982 18860 31034
rect 1104 30960 18860 30982
rect 6454 30812 6460 30864
rect 6512 30812 6518 30864
rect 5718 30744 5724 30796
rect 5776 30784 5782 30796
rect 6472 30784 6500 30812
rect 5776 30756 6132 30784
rect 6472 30756 8064 30784
rect 5776 30744 5782 30756
rect 934 30676 940 30728
rect 992 30716 998 30728
rect 1581 30719 1639 30725
rect 1581 30716 1593 30719
rect 992 30688 1593 30716
rect 992 30676 998 30688
rect 1581 30685 1593 30688
rect 1627 30685 1639 30719
rect 1581 30679 1639 30685
rect 5994 30676 6000 30728
rect 6052 30676 6058 30728
rect 6104 30725 6132 30756
rect 6089 30719 6147 30725
rect 6089 30685 6101 30719
rect 6135 30685 6147 30719
rect 6089 30679 6147 30685
rect 6362 30676 6368 30728
rect 6420 30716 6426 30728
rect 6457 30719 6515 30725
rect 6457 30716 6469 30719
rect 6420 30688 6469 30716
rect 6420 30676 6426 30688
rect 6457 30685 6469 30688
rect 6503 30716 6515 30719
rect 7101 30719 7159 30725
rect 6503 30688 6868 30716
rect 6503 30685 6515 30688
rect 6457 30679 6515 30685
rect 5721 30651 5779 30657
rect 5721 30617 5733 30651
rect 5767 30648 5779 30651
rect 6546 30648 6552 30660
rect 5767 30620 6552 30648
rect 5767 30617 5779 30620
rect 5721 30611 5779 30617
rect 6546 30608 6552 30620
rect 6604 30608 6610 30660
rect 6840 30648 6868 30688
rect 7101 30685 7113 30719
rect 7147 30716 7159 30719
rect 7147 30688 7420 30716
rect 7147 30685 7159 30688
rect 7101 30679 7159 30685
rect 7190 30648 7196 30660
rect 6840 30620 7196 30648
rect 7190 30608 7196 30620
rect 7248 30608 7254 30660
rect 7392 30648 7420 30688
rect 7466 30676 7472 30728
rect 7524 30676 7530 30728
rect 8036 30725 8064 30756
rect 8021 30719 8079 30725
rect 8021 30685 8033 30719
rect 8067 30685 8079 30719
rect 8021 30679 8079 30685
rect 7558 30648 7564 30660
rect 7392 30620 7564 30648
rect 7558 30608 7564 30620
rect 7616 30608 7622 30660
rect 5994 30540 6000 30592
rect 6052 30580 6058 30592
rect 6914 30580 6920 30592
rect 6052 30552 6920 30580
rect 6052 30540 6058 30552
rect 6914 30540 6920 30552
rect 6972 30540 6978 30592
rect 8018 30540 8024 30592
rect 8076 30580 8082 30592
rect 8205 30583 8263 30589
rect 8205 30580 8217 30583
rect 8076 30552 8217 30580
rect 8076 30540 8082 30552
rect 8205 30549 8217 30552
rect 8251 30549 8263 30583
rect 8205 30543 8263 30549
rect 1104 30490 19019 30512
rect 1104 30438 5388 30490
rect 5440 30438 5452 30490
rect 5504 30438 5516 30490
rect 5568 30438 5580 30490
rect 5632 30438 5644 30490
rect 5696 30438 9827 30490
rect 9879 30438 9891 30490
rect 9943 30438 9955 30490
rect 10007 30438 10019 30490
rect 10071 30438 10083 30490
rect 10135 30438 14266 30490
rect 14318 30438 14330 30490
rect 14382 30438 14394 30490
rect 14446 30438 14458 30490
rect 14510 30438 14522 30490
rect 14574 30438 18705 30490
rect 18757 30438 18769 30490
rect 18821 30438 18833 30490
rect 18885 30438 18897 30490
rect 18949 30438 18961 30490
rect 19013 30438 19019 30490
rect 1104 30416 19019 30438
rect 6730 30336 6736 30388
rect 6788 30376 6794 30388
rect 7558 30376 7564 30388
rect 6788 30348 7564 30376
rect 6788 30336 6794 30348
rect 7558 30336 7564 30348
rect 7616 30376 7622 30388
rect 8938 30376 8944 30388
rect 7616 30348 8944 30376
rect 7616 30336 7622 30348
rect 8938 30336 8944 30348
rect 8996 30336 9002 30388
rect 6178 30268 6184 30320
rect 6236 30308 6242 30320
rect 6236 30280 7328 30308
rect 6236 30268 6242 30280
rect 7006 30200 7012 30252
rect 7064 30200 7070 30252
rect 7300 30249 7328 30280
rect 7285 30243 7343 30249
rect 7285 30209 7297 30243
rect 7331 30209 7343 30243
rect 7285 30203 7343 30209
rect 7469 30243 7527 30249
rect 7469 30209 7481 30243
rect 7515 30240 7527 30243
rect 7926 30240 7932 30252
rect 7515 30212 7932 30240
rect 7515 30209 7527 30212
rect 7469 30203 7527 30209
rect 7190 30132 7196 30184
rect 7248 30172 7254 30184
rect 7484 30172 7512 30203
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 8021 30243 8079 30249
rect 8021 30209 8033 30243
rect 8067 30209 8079 30243
rect 8021 30203 8079 30209
rect 8036 30172 8064 30203
rect 7248 30144 7512 30172
rect 7944 30144 8064 30172
rect 7248 30132 7254 30144
rect 7374 30064 7380 30116
rect 7432 30064 7438 30116
rect 6822 29996 6828 30048
rect 6880 30036 6886 30048
rect 7944 30036 7972 30144
rect 6880 30008 7972 30036
rect 6880 29996 6886 30008
rect 8110 29996 8116 30048
rect 8168 29996 8174 30048
rect 1104 29946 18860 29968
rect 1104 29894 3169 29946
rect 3221 29894 3233 29946
rect 3285 29894 3297 29946
rect 3349 29894 3361 29946
rect 3413 29894 3425 29946
rect 3477 29894 7608 29946
rect 7660 29894 7672 29946
rect 7724 29894 7736 29946
rect 7788 29894 7800 29946
rect 7852 29894 7864 29946
rect 7916 29894 12047 29946
rect 12099 29894 12111 29946
rect 12163 29894 12175 29946
rect 12227 29894 12239 29946
rect 12291 29894 12303 29946
rect 12355 29894 16486 29946
rect 16538 29894 16550 29946
rect 16602 29894 16614 29946
rect 16666 29894 16678 29946
rect 16730 29894 16742 29946
rect 16794 29894 18860 29946
rect 1104 29872 18860 29894
rect 5629 29835 5687 29841
rect 5629 29801 5641 29835
rect 5675 29832 5687 29835
rect 5718 29832 5724 29844
rect 5675 29804 5724 29832
rect 5675 29801 5687 29804
rect 5629 29795 5687 29801
rect 5718 29792 5724 29804
rect 5776 29792 5782 29844
rect 7466 29792 7472 29844
rect 7524 29792 7530 29844
rect 7006 29724 7012 29776
rect 7064 29764 7070 29776
rect 8202 29764 8208 29776
rect 7064 29736 8208 29764
rect 7064 29724 7070 29736
rect 8202 29724 8208 29736
rect 8260 29724 8266 29776
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29628 4951 29631
rect 4982 29628 4988 29640
rect 4939 29600 4988 29628
rect 4939 29597 4951 29600
rect 4893 29591 4951 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 6178 29588 6184 29640
rect 6236 29588 6242 29640
rect 6730 29588 6736 29640
rect 6788 29588 6794 29640
rect 6917 29631 6975 29637
rect 6917 29597 6929 29631
rect 6963 29628 6975 29631
rect 7006 29628 7012 29640
rect 6963 29600 7012 29628
rect 6963 29597 6975 29600
rect 6917 29591 6975 29597
rect 7006 29588 7012 29600
rect 7064 29588 7070 29640
rect 7374 29588 7380 29640
rect 7432 29628 7438 29640
rect 7561 29631 7619 29637
rect 7561 29628 7573 29631
rect 7432 29600 7573 29628
rect 7432 29588 7438 29600
rect 7561 29597 7573 29600
rect 7607 29597 7619 29631
rect 7561 29591 7619 29597
rect 5074 29520 5080 29572
rect 5132 29560 5138 29572
rect 5169 29563 5227 29569
rect 5169 29560 5181 29563
rect 5132 29532 5181 29560
rect 5132 29520 5138 29532
rect 5169 29529 5181 29532
rect 5215 29529 5227 29563
rect 5169 29523 5227 29529
rect 4614 29452 4620 29504
rect 4672 29452 4678 29504
rect 4798 29452 4804 29504
rect 4856 29452 4862 29504
rect 4890 29452 4896 29504
rect 4948 29492 4954 29504
rect 4985 29495 5043 29501
rect 4985 29492 4997 29495
rect 4948 29464 4997 29492
rect 4948 29452 4954 29464
rect 4985 29461 4997 29464
rect 5031 29461 5043 29495
rect 4985 29455 5043 29461
rect 1104 29402 19019 29424
rect 1104 29350 5388 29402
rect 5440 29350 5452 29402
rect 5504 29350 5516 29402
rect 5568 29350 5580 29402
rect 5632 29350 5644 29402
rect 5696 29350 9827 29402
rect 9879 29350 9891 29402
rect 9943 29350 9955 29402
rect 10007 29350 10019 29402
rect 10071 29350 10083 29402
rect 10135 29350 14266 29402
rect 14318 29350 14330 29402
rect 14382 29350 14394 29402
rect 14446 29350 14458 29402
rect 14510 29350 14522 29402
rect 14574 29350 18705 29402
rect 18757 29350 18769 29402
rect 18821 29350 18833 29402
rect 18885 29350 18897 29402
rect 18949 29350 18961 29402
rect 19013 29350 19019 29402
rect 1104 29328 19019 29350
rect 6914 29248 6920 29300
rect 6972 29248 6978 29300
rect 7466 29248 7472 29300
rect 7524 29288 7530 29300
rect 7929 29291 7987 29297
rect 7929 29288 7941 29291
rect 7524 29260 7941 29288
rect 7524 29248 7530 29260
rect 7929 29257 7941 29260
rect 7975 29257 7987 29291
rect 7929 29251 7987 29257
rect 4890 29180 4896 29232
rect 4948 29180 4954 29232
rect 6932 29220 6960 29248
rect 6932 29192 7512 29220
rect 4522 29112 4528 29164
rect 4580 29152 4586 29164
rect 4908 29152 4936 29180
rect 7484 29164 7512 29192
rect 5169 29155 5227 29161
rect 5169 29152 5181 29155
rect 4580 29124 5181 29152
rect 4580 29112 4586 29124
rect 5169 29121 5181 29124
rect 5215 29121 5227 29155
rect 5169 29115 5227 29121
rect 6549 29155 6607 29161
rect 6549 29121 6561 29155
rect 6595 29121 6607 29155
rect 6549 29115 6607 29121
rect 4798 29044 4804 29096
rect 4856 29084 4862 29096
rect 4893 29087 4951 29093
rect 4893 29084 4905 29087
rect 4856 29056 4905 29084
rect 4856 29044 4862 29056
rect 4893 29053 4905 29056
rect 4939 29053 4951 29087
rect 4893 29047 4951 29053
rect 4982 29044 4988 29096
rect 5040 29044 5046 29096
rect 5074 29044 5080 29096
rect 5132 29044 5138 29096
rect 6564 29084 6592 29115
rect 6638 29112 6644 29164
rect 6696 29112 6702 29164
rect 6822 29112 6828 29164
rect 6880 29112 6886 29164
rect 6917 29155 6975 29161
rect 6917 29121 6929 29155
rect 6963 29152 6975 29155
rect 7098 29152 7104 29164
rect 6963 29124 7104 29152
rect 6963 29121 6975 29124
rect 6917 29115 6975 29121
rect 7098 29112 7104 29124
rect 7156 29112 7162 29164
rect 7466 29112 7472 29164
rect 7524 29152 7530 29164
rect 7745 29155 7803 29161
rect 7745 29152 7757 29155
rect 7524 29124 7757 29152
rect 7524 29112 7530 29124
rect 7745 29121 7757 29124
rect 7791 29121 7803 29155
rect 7745 29115 7803 29121
rect 8018 29112 8024 29164
rect 8076 29112 8082 29164
rect 6730 29084 6736 29096
rect 6564 29056 6736 29084
rect 6730 29044 6736 29056
rect 6788 29044 6794 29096
rect 6454 28976 6460 29028
rect 6512 29016 6518 29028
rect 7561 29019 7619 29025
rect 7561 29016 7573 29019
rect 6512 28988 7573 29016
rect 6512 28976 6518 28988
rect 7561 28985 7573 28988
rect 7607 28985 7619 29019
rect 7561 28979 7619 28985
rect 4706 28908 4712 28960
rect 4764 28908 4770 28960
rect 5258 28908 5264 28960
rect 5316 28948 5322 28960
rect 7101 28951 7159 28957
rect 7101 28948 7113 28951
rect 5316 28920 7113 28948
rect 5316 28908 5322 28920
rect 7101 28917 7113 28920
rect 7147 28917 7159 28951
rect 7101 28911 7159 28917
rect 1104 28858 18860 28880
rect 1104 28806 3169 28858
rect 3221 28806 3233 28858
rect 3285 28806 3297 28858
rect 3349 28806 3361 28858
rect 3413 28806 3425 28858
rect 3477 28806 7608 28858
rect 7660 28806 7672 28858
rect 7724 28806 7736 28858
rect 7788 28806 7800 28858
rect 7852 28806 7864 28858
rect 7916 28806 12047 28858
rect 12099 28806 12111 28858
rect 12163 28806 12175 28858
rect 12227 28806 12239 28858
rect 12291 28806 12303 28858
rect 12355 28806 16486 28858
rect 16538 28806 16550 28858
rect 16602 28806 16614 28858
rect 16666 28806 16678 28858
rect 16730 28806 16742 28858
rect 16794 28806 18860 28858
rect 1104 28784 18860 28806
rect 4154 28704 4160 28756
rect 4212 28744 4218 28756
rect 4433 28747 4491 28753
rect 4433 28744 4445 28747
rect 4212 28716 4445 28744
rect 4212 28704 4218 28716
rect 4433 28713 4445 28716
rect 4479 28713 4491 28747
rect 4433 28707 4491 28713
rect 4614 28636 4620 28688
rect 4672 28676 4678 28688
rect 4801 28679 4859 28685
rect 4801 28676 4813 28679
rect 4672 28648 4813 28676
rect 4672 28636 4678 28648
rect 4801 28645 4813 28648
rect 4847 28676 4859 28679
rect 5718 28676 5724 28688
rect 4847 28648 5724 28676
rect 4847 28645 4859 28648
rect 4801 28639 4859 28645
rect 5718 28636 5724 28648
rect 5776 28636 5782 28688
rect 6454 28568 6460 28620
rect 6512 28568 6518 28620
rect 6641 28611 6699 28617
rect 6641 28577 6653 28611
rect 6687 28608 6699 28611
rect 6822 28608 6828 28620
rect 6687 28580 6828 28608
rect 6687 28577 6699 28580
rect 6641 28571 6699 28577
rect 6822 28568 6828 28580
rect 6880 28608 6886 28620
rect 8021 28611 8079 28617
rect 8021 28608 8033 28611
rect 6880 28580 8033 28608
rect 6880 28568 6886 28580
rect 8021 28577 8033 28580
rect 8067 28577 8079 28611
rect 8021 28571 8079 28577
rect 3237 28543 3295 28549
rect 3237 28509 3249 28543
rect 3283 28509 3295 28543
rect 3237 28503 3295 28509
rect 3421 28543 3479 28549
rect 3421 28509 3433 28543
rect 3467 28540 3479 28543
rect 4062 28540 4068 28552
rect 3467 28512 4068 28540
rect 3467 28509 3479 28512
rect 3421 28503 3479 28509
rect 3252 28472 3280 28503
rect 4062 28500 4068 28512
rect 4120 28500 4126 28552
rect 6546 28500 6552 28552
rect 6604 28500 6610 28552
rect 6730 28500 6736 28552
rect 6788 28540 6794 28552
rect 7282 28540 7288 28552
rect 6788 28512 7288 28540
rect 6788 28500 6794 28512
rect 7282 28500 7288 28512
rect 7340 28500 7346 28552
rect 7466 28500 7472 28552
rect 7524 28500 7530 28552
rect 7653 28543 7711 28549
rect 7653 28509 7665 28543
rect 7699 28540 7711 28543
rect 7926 28540 7932 28552
rect 7699 28512 7932 28540
rect 7699 28509 7711 28512
rect 7653 28503 7711 28509
rect 7926 28500 7932 28512
rect 7984 28500 7990 28552
rect 3786 28472 3792 28484
rect 3252 28444 3792 28472
rect 3786 28432 3792 28444
rect 3844 28432 3850 28484
rect 4433 28475 4491 28481
rect 4433 28441 4445 28475
rect 4479 28472 4491 28475
rect 4706 28472 4712 28484
rect 4479 28444 4712 28472
rect 4479 28441 4491 28444
rect 4433 28435 4491 28441
rect 4706 28432 4712 28444
rect 4764 28432 4770 28484
rect 3329 28407 3387 28413
rect 3329 28373 3341 28407
rect 3375 28404 3387 28407
rect 3970 28404 3976 28416
rect 3375 28376 3976 28404
rect 3375 28373 3387 28376
rect 3329 28367 3387 28373
rect 3970 28364 3976 28376
rect 4028 28364 4034 28416
rect 4246 28364 4252 28416
rect 4304 28364 4310 28416
rect 6270 28364 6276 28416
rect 6328 28364 6334 28416
rect 7282 28364 7288 28416
rect 7340 28404 7346 28416
rect 7929 28407 7987 28413
rect 7929 28404 7941 28407
rect 7340 28376 7941 28404
rect 7340 28364 7346 28376
rect 7929 28373 7941 28376
rect 7975 28373 7987 28407
rect 7929 28367 7987 28373
rect 1104 28314 19019 28336
rect 1104 28262 5388 28314
rect 5440 28262 5452 28314
rect 5504 28262 5516 28314
rect 5568 28262 5580 28314
rect 5632 28262 5644 28314
rect 5696 28262 9827 28314
rect 9879 28262 9891 28314
rect 9943 28262 9955 28314
rect 10007 28262 10019 28314
rect 10071 28262 10083 28314
rect 10135 28262 14266 28314
rect 14318 28262 14330 28314
rect 14382 28262 14394 28314
rect 14446 28262 14458 28314
rect 14510 28262 14522 28314
rect 14574 28262 18705 28314
rect 18757 28262 18769 28314
rect 18821 28262 18833 28314
rect 18885 28262 18897 28314
rect 18949 28262 18961 28314
rect 19013 28262 19019 28314
rect 1104 28240 19019 28262
rect 6454 28024 6460 28076
rect 6512 28064 6518 28076
rect 8573 28067 8631 28073
rect 8573 28064 8585 28067
rect 6512 28036 8585 28064
rect 6512 28024 6518 28036
rect 8573 28033 8585 28036
rect 8619 28033 8631 28067
rect 8573 28027 8631 28033
rect 8849 28067 8907 28073
rect 8849 28033 8861 28067
rect 8895 28064 8907 28067
rect 8938 28064 8944 28076
rect 8895 28036 8944 28064
rect 8895 28033 8907 28036
rect 8849 28027 8907 28033
rect 8938 28024 8944 28036
rect 8996 28024 9002 28076
rect 8018 27956 8024 28008
rect 8076 27996 8082 28008
rect 8481 27999 8539 28005
rect 8481 27996 8493 27999
rect 8076 27968 8493 27996
rect 8076 27956 8082 27968
rect 8481 27965 8493 27968
rect 8527 27965 8539 27999
rect 8481 27959 8539 27965
rect 1104 27770 18860 27792
rect 1104 27718 3169 27770
rect 3221 27718 3233 27770
rect 3285 27718 3297 27770
rect 3349 27718 3361 27770
rect 3413 27718 3425 27770
rect 3477 27718 7608 27770
rect 7660 27718 7672 27770
rect 7724 27718 7736 27770
rect 7788 27718 7800 27770
rect 7852 27718 7864 27770
rect 7916 27718 12047 27770
rect 12099 27718 12111 27770
rect 12163 27718 12175 27770
rect 12227 27718 12239 27770
rect 12291 27718 12303 27770
rect 12355 27718 16486 27770
rect 16538 27718 16550 27770
rect 16602 27718 16614 27770
rect 16666 27718 16678 27770
rect 16730 27718 16742 27770
rect 16794 27718 18860 27770
rect 1104 27696 18860 27718
rect 3329 27591 3387 27597
rect 3329 27557 3341 27591
rect 3375 27588 3387 27591
rect 4246 27588 4252 27600
rect 3375 27560 4252 27588
rect 3375 27557 3387 27560
rect 3329 27551 3387 27557
rect 4246 27548 4252 27560
rect 4304 27548 4310 27600
rect 3421 27523 3479 27529
rect 3421 27489 3433 27523
rect 3467 27520 3479 27523
rect 3602 27520 3608 27532
rect 3467 27492 3608 27520
rect 3467 27489 3479 27492
rect 3421 27483 3479 27489
rect 3602 27480 3608 27492
rect 3660 27480 3666 27532
rect 5810 27520 5816 27532
rect 3712 27492 5816 27520
rect 3145 27455 3203 27461
rect 3145 27421 3157 27455
rect 3191 27421 3203 27455
rect 3145 27415 3203 27421
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27452 3295 27455
rect 3712 27452 3740 27492
rect 5810 27480 5816 27492
rect 5868 27480 5874 27532
rect 3283 27424 3740 27452
rect 3283 27421 3295 27424
rect 3237 27415 3295 27421
rect 3160 27316 3188 27415
rect 3786 27412 3792 27464
rect 3844 27452 3850 27464
rect 3973 27455 4031 27461
rect 3973 27452 3985 27455
rect 3844 27424 3985 27452
rect 3844 27412 3850 27424
rect 3973 27421 3985 27424
rect 4019 27421 4031 27455
rect 3973 27415 4031 27421
rect 4062 27412 4068 27464
rect 4120 27452 4126 27464
rect 4249 27455 4307 27461
rect 4249 27452 4261 27455
rect 4120 27424 4261 27452
rect 4120 27412 4126 27424
rect 4249 27421 4261 27424
rect 4295 27421 4307 27455
rect 4249 27415 4307 27421
rect 4430 27412 4436 27464
rect 4488 27412 4494 27464
rect 4614 27412 4620 27464
rect 4672 27412 4678 27464
rect 4801 27387 4859 27393
rect 4801 27353 4813 27387
rect 4847 27384 4859 27387
rect 6822 27384 6828 27396
rect 4847 27356 6828 27384
rect 4847 27353 4859 27356
rect 4801 27347 4859 27353
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 6638 27316 6644 27328
rect 3160 27288 6644 27316
rect 6638 27276 6644 27288
rect 6696 27276 6702 27328
rect 1104 27226 19019 27248
rect 1104 27174 5388 27226
rect 5440 27174 5452 27226
rect 5504 27174 5516 27226
rect 5568 27174 5580 27226
rect 5632 27174 5644 27226
rect 5696 27174 9827 27226
rect 9879 27174 9891 27226
rect 9943 27174 9955 27226
rect 10007 27174 10019 27226
rect 10071 27174 10083 27226
rect 10135 27174 14266 27226
rect 14318 27174 14330 27226
rect 14382 27174 14394 27226
rect 14446 27174 14458 27226
rect 14510 27174 14522 27226
rect 14574 27174 18705 27226
rect 18757 27174 18769 27226
rect 18821 27174 18833 27226
rect 18885 27174 18897 27226
rect 18949 27174 18961 27226
rect 19013 27174 19019 27226
rect 1104 27152 19019 27174
rect 3602 27072 3608 27124
rect 3660 27112 3666 27124
rect 4154 27112 4160 27124
rect 3660 27084 4160 27112
rect 3660 27072 3666 27084
rect 4154 27072 4160 27084
rect 4212 27072 4218 27124
rect 4617 27115 4675 27121
rect 4617 27081 4629 27115
rect 4663 27112 4675 27115
rect 4982 27112 4988 27124
rect 4663 27084 4988 27112
rect 4663 27081 4675 27084
rect 4617 27075 4675 27081
rect 4982 27072 4988 27084
rect 5040 27072 5046 27124
rect 2866 27004 2872 27056
rect 2924 27044 2930 27056
rect 4062 27044 4068 27056
rect 2924 27016 4068 27044
rect 2924 27004 2930 27016
rect 4062 27004 4068 27016
rect 4120 27004 4126 27056
rect 6178 27004 6184 27056
rect 6236 27044 6242 27056
rect 6549 27047 6607 27053
rect 6549 27044 6561 27047
rect 6236 27016 6561 27044
rect 6236 27004 6242 27016
rect 6549 27013 6561 27016
rect 6595 27013 6607 27047
rect 6549 27007 6607 27013
rect 6822 27004 6828 27056
rect 6880 27044 6886 27056
rect 6917 27047 6975 27053
rect 6917 27044 6929 27047
rect 6880 27016 6929 27044
rect 6880 27004 6886 27016
rect 6917 27013 6929 27016
rect 6963 27013 6975 27047
rect 6917 27007 6975 27013
rect 7009 27047 7067 27053
rect 7009 27013 7021 27047
rect 7055 27044 7067 27047
rect 7466 27044 7472 27056
rect 7055 27016 7472 27044
rect 7055 27013 7067 27016
rect 7009 27007 7067 27013
rect 7466 27004 7472 27016
rect 7524 27004 7530 27056
rect 1762 26936 1768 26988
rect 1820 26936 1826 26988
rect 4338 26936 4344 26988
rect 4396 26976 4402 26988
rect 4433 26979 4491 26985
rect 4433 26976 4445 26979
rect 4396 26948 4445 26976
rect 4396 26936 4402 26948
rect 4433 26945 4445 26948
rect 4479 26945 4491 26979
rect 4433 26939 4491 26945
rect 5626 26936 5632 26988
rect 5684 26936 5690 26988
rect 5721 26979 5779 26985
rect 5721 26945 5733 26979
rect 5767 26976 5779 26979
rect 6362 26976 6368 26988
rect 5767 26948 6368 26976
rect 5767 26945 5779 26948
rect 5721 26939 5779 26945
rect 6362 26936 6368 26948
rect 6420 26936 6426 26988
rect 7101 26979 7159 26985
rect 7101 26945 7113 26979
rect 7147 26945 7159 26979
rect 7101 26939 7159 26945
rect 2130 26868 2136 26920
rect 2188 26908 2194 26920
rect 4249 26911 4307 26917
rect 4249 26908 4261 26911
rect 2188 26880 4261 26908
rect 2188 26868 2194 26880
rect 4249 26877 4261 26880
rect 4295 26908 4307 26911
rect 4890 26908 4896 26920
rect 4295 26880 4896 26908
rect 4295 26877 4307 26880
rect 4249 26871 4307 26877
rect 4890 26868 4896 26880
rect 4948 26868 4954 26920
rect 6914 26868 6920 26920
rect 6972 26908 6978 26920
rect 7116 26908 7144 26939
rect 6972 26880 7144 26908
rect 7285 26911 7343 26917
rect 6972 26868 6978 26880
rect 7285 26877 7297 26911
rect 7331 26908 7343 26911
rect 7374 26908 7380 26920
rect 7331 26880 7380 26908
rect 7331 26877 7343 26880
rect 7285 26871 7343 26877
rect 7374 26868 7380 26880
rect 7432 26868 7438 26920
rect 8021 26911 8079 26917
rect 8021 26877 8033 26911
rect 8067 26877 8079 26911
rect 8021 26871 8079 26877
rect 934 26800 940 26852
rect 992 26840 998 26852
rect 1581 26843 1639 26849
rect 1581 26840 1593 26843
rect 992 26812 1593 26840
rect 992 26800 998 26812
rect 1581 26809 1593 26812
rect 1627 26809 1639 26843
rect 1581 26803 1639 26809
rect 6730 26800 6736 26852
rect 6788 26840 6794 26852
rect 8036 26840 8064 26871
rect 6788 26812 8064 26840
rect 6788 26800 6794 26812
rect 8294 26800 8300 26852
rect 8352 26800 8358 26852
rect 5902 26732 5908 26784
rect 5960 26732 5966 26784
rect 8478 26732 8484 26784
rect 8536 26732 8542 26784
rect 1104 26682 18860 26704
rect 1104 26630 3169 26682
rect 3221 26630 3233 26682
rect 3285 26630 3297 26682
rect 3349 26630 3361 26682
rect 3413 26630 3425 26682
rect 3477 26630 7608 26682
rect 7660 26630 7672 26682
rect 7724 26630 7736 26682
rect 7788 26630 7800 26682
rect 7852 26630 7864 26682
rect 7916 26630 12047 26682
rect 12099 26630 12111 26682
rect 12163 26630 12175 26682
rect 12227 26630 12239 26682
rect 12291 26630 12303 26682
rect 12355 26630 16486 26682
rect 16538 26630 16550 26682
rect 16602 26630 16614 26682
rect 16666 26630 16678 26682
rect 16730 26630 16742 26682
rect 16794 26630 18860 26682
rect 1104 26608 18860 26630
rect 4341 26571 4399 26577
rect 4341 26537 4353 26571
rect 4387 26568 4399 26571
rect 4430 26568 4436 26580
rect 4387 26540 4436 26568
rect 4387 26537 4399 26540
rect 4341 26531 4399 26537
rect 4430 26528 4436 26540
rect 4488 26528 4494 26580
rect 4522 26528 4528 26580
rect 4580 26528 4586 26580
rect 4706 26460 4712 26512
rect 4764 26500 4770 26512
rect 6270 26500 6276 26512
rect 4764 26472 6276 26500
rect 4764 26460 4770 26472
rect 6270 26460 6276 26472
rect 6328 26460 6334 26512
rect 6641 26503 6699 26509
rect 6641 26469 6653 26503
rect 6687 26500 6699 26503
rect 8754 26500 8760 26512
rect 6687 26472 8760 26500
rect 6687 26469 6699 26472
rect 6641 26463 6699 26469
rect 8754 26460 8760 26472
rect 8812 26460 8818 26512
rect 2590 26392 2596 26444
rect 2648 26432 2654 26444
rect 4338 26432 4344 26444
rect 2648 26404 4344 26432
rect 2648 26392 2654 26404
rect 4338 26392 4344 26404
rect 4396 26432 4402 26444
rect 4985 26435 5043 26441
rect 4985 26432 4997 26435
rect 4396 26404 4997 26432
rect 4396 26392 4402 26404
rect 4985 26401 4997 26404
rect 5031 26401 5043 26435
rect 4985 26395 5043 26401
rect 6086 26392 6092 26444
rect 6144 26432 6150 26444
rect 7009 26435 7067 26441
rect 7009 26432 7021 26435
rect 6144 26404 7021 26432
rect 6144 26392 6150 26404
rect 7009 26401 7021 26404
rect 7055 26401 7067 26435
rect 7009 26395 7067 26401
rect 4525 26367 4583 26373
rect 4525 26333 4537 26367
rect 4571 26333 4583 26367
rect 4525 26327 4583 26333
rect 4540 26296 4568 26327
rect 4890 26324 4896 26376
rect 4948 26324 4954 26376
rect 5810 26324 5816 26376
rect 5868 26324 5874 26376
rect 5994 26324 6000 26376
rect 6052 26324 6058 26376
rect 6454 26324 6460 26376
rect 6512 26364 6518 26376
rect 6825 26367 6883 26373
rect 6825 26364 6837 26367
rect 6512 26336 6837 26364
rect 6512 26324 6518 26336
rect 6825 26333 6837 26336
rect 6871 26333 6883 26367
rect 6825 26327 6883 26333
rect 6917 26367 6975 26373
rect 6917 26333 6929 26367
rect 6963 26333 6975 26367
rect 6917 26327 6975 26333
rect 7101 26367 7159 26373
rect 7101 26333 7113 26367
rect 7147 26364 7159 26367
rect 7282 26364 7288 26376
rect 7147 26336 7288 26364
rect 7147 26333 7159 26336
rect 7101 26327 7159 26333
rect 5074 26296 5080 26308
rect 4540 26268 5080 26296
rect 2038 26188 2044 26240
rect 2096 26228 2102 26240
rect 4540 26228 4568 26268
rect 5074 26256 5080 26268
rect 5132 26256 5138 26308
rect 6178 26256 6184 26308
rect 6236 26256 6242 26308
rect 6932 26296 6960 26327
rect 7282 26324 7288 26336
rect 7340 26324 7346 26376
rect 7926 26296 7932 26308
rect 6932 26268 7932 26296
rect 7926 26256 7932 26268
rect 7984 26296 7990 26308
rect 8570 26296 8576 26308
rect 7984 26268 8576 26296
rect 7984 26256 7990 26268
rect 8570 26256 8576 26268
rect 8628 26256 8634 26308
rect 2096 26200 4568 26228
rect 2096 26188 2102 26200
rect 8202 26188 8208 26240
rect 8260 26228 8266 26240
rect 8386 26228 8392 26240
rect 8260 26200 8392 26228
rect 8260 26188 8266 26200
rect 8386 26188 8392 26200
rect 8444 26188 8450 26240
rect 1104 26138 19019 26160
rect 1104 26086 5388 26138
rect 5440 26086 5452 26138
rect 5504 26086 5516 26138
rect 5568 26086 5580 26138
rect 5632 26086 5644 26138
rect 5696 26086 9827 26138
rect 9879 26086 9891 26138
rect 9943 26086 9955 26138
rect 10007 26086 10019 26138
rect 10071 26086 10083 26138
rect 10135 26086 14266 26138
rect 14318 26086 14330 26138
rect 14382 26086 14394 26138
rect 14446 26086 14458 26138
rect 14510 26086 14522 26138
rect 14574 26086 18705 26138
rect 18757 26086 18769 26138
rect 18821 26086 18833 26138
rect 18885 26086 18897 26138
rect 18949 26086 18961 26138
rect 19013 26086 19019 26138
rect 1104 26064 19019 26086
rect 6549 26027 6607 26033
rect 6549 25993 6561 26027
rect 6595 26024 6607 26027
rect 7006 26024 7012 26036
rect 6595 25996 7012 26024
rect 6595 25993 6607 25996
rect 6549 25987 6607 25993
rect 7006 25984 7012 25996
rect 7064 25984 7070 26036
rect 4430 25956 4436 25968
rect 3988 25928 4436 25956
rect 3988 25897 4016 25928
rect 4430 25916 4436 25928
rect 4488 25916 4494 25968
rect 6822 25956 6828 25968
rect 6748 25928 6828 25956
rect 3973 25891 4031 25897
rect 3973 25857 3985 25891
rect 4019 25857 4031 25891
rect 3973 25851 4031 25857
rect 4157 25891 4215 25897
rect 4157 25857 4169 25891
rect 4203 25888 4215 25891
rect 4338 25888 4344 25900
rect 4203 25860 4344 25888
rect 4203 25857 4215 25860
rect 4157 25851 4215 25857
rect 4338 25848 4344 25860
rect 4396 25888 4402 25900
rect 4614 25888 4620 25900
rect 4396 25860 4620 25888
rect 4396 25848 4402 25860
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 6748 25897 6776 25928
rect 6822 25916 6828 25928
rect 6880 25916 6886 25968
rect 6733 25891 6791 25897
rect 6733 25857 6745 25891
rect 6779 25857 6791 25891
rect 7466 25888 7472 25900
rect 6733 25851 6791 25857
rect 6840 25860 7472 25888
rect 5074 25780 5080 25832
rect 5132 25820 5138 25832
rect 6840 25829 6868 25860
rect 7466 25848 7472 25860
rect 7524 25848 7530 25900
rect 6825 25823 6883 25829
rect 6825 25820 6837 25823
rect 5132 25792 6837 25820
rect 5132 25780 5138 25792
rect 6825 25789 6837 25792
rect 6871 25789 6883 25823
rect 6825 25783 6883 25789
rect 6914 25780 6920 25832
rect 6972 25780 6978 25832
rect 7009 25823 7067 25829
rect 7009 25789 7021 25823
rect 7055 25820 7067 25823
rect 7374 25820 7380 25832
rect 7055 25792 7380 25820
rect 7055 25789 7067 25792
rect 7009 25783 7067 25789
rect 7374 25780 7380 25792
rect 7432 25780 7438 25832
rect 4157 25687 4215 25693
rect 4157 25653 4169 25687
rect 4203 25684 4215 25687
rect 5166 25684 5172 25696
rect 4203 25656 5172 25684
rect 4203 25653 4215 25656
rect 4157 25647 4215 25653
rect 5166 25644 5172 25656
rect 5224 25644 5230 25696
rect 1104 25594 18860 25616
rect 1104 25542 3169 25594
rect 3221 25542 3233 25594
rect 3285 25542 3297 25594
rect 3349 25542 3361 25594
rect 3413 25542 3425 25594
rect 3477 25542 7608 25594
rect 7660 25542 7672 25594
rect 7724 25542 7736 25594
rect 7788 25542 7800 25594
rect 7852 25542 7864 25594
rect 7916 25542 12047 25594
rect 12099 25542 12111 25594
rect 12163 25542 12175 25594
rect 12227 25542 12239 25594
rect 12291 25542 12303 25594
rect 12355 25542 16486 25594
rect 16538 25542 16550 25594
rect 16602 25542 16614 25594
rect 16666 25542 16678 25594
rect 16730 25542 16742 25594
rect 16794 25542 18860 25594
rect 1104 25520 18860 25542
rect 2130 25440 2136 25492
rect 2188 25440 2194 25492
rect 5810 25440 5816 25492
rect 5868 25480 5874 25492
rect 6273 25483 6331 25489
rect 6273 25480 6285 25483
rect 5868 25452 6285 25480
rect 5868 25440 5874 25452
rect 6273 25449 6285 25452
rect 6319 25449 6331 25483
rect 6273 25443 6331 25449
rect 6457 25483 6515 25489
rect 6457 25449 6469 25483
rect 6503 25449 6515 25483
rect 6457 25443 6515 25449
rect 5718 25372 5724 25424
rect 5776 25412 5782 25424
rect 6472 25412 6500 25443
rect 8110 25440 8116 25492
rect 8168 25440 8174 25492
rect 5776 25384 6500 25412
rect 5776 25372 5782 25384
rect 5537 25347 5595 25353
rect 5537 25313 5549 25347
rect 5583 25344 5595 25347
rect 7006 25344 7012 25356
rect 5583 25316 7012 25344
rect 5583 25313 5595 25316
rect 5537 25307 5595 25313
rect 7006 25304 7012 25316
rect 7064 25304 7070 25356
rect 3602 25236 3608 25288
rect 3660 25276 3666 25288
rect 4062 25276 4068 25288
rect 3660 25248 4068 25276
rect 3660 25236 3666 25248
rect 4062 25236 4068 25248
rect 4120 25276 4126 25288
rect 5353 25279 5411 25285
rect 5353 25276 5365 25279
rect 4120 25248 5365 25276
rect 4120 25236 4126 25248
rect 5353 25245 5365 25248
rect 5399 25245 5411 25279
rect 5353 25239 5411 25245
rect 5810 25236 5816 25288
rect 5868 25236 5874 25288
rect 7834 25236 7840 25288
rect 7892 25236 7898 25288
rect 2038 25168 2044 25220
rect 2096 25208 2102 25220
rect 2317 25211 2375 25217
rect 2317 25208 2329 25211
rect 2096 25180 2329 25208
rect 2096 25168 2102 25180
rect 2317 25177 2329 25180
rect 2363 25177 2375 25211
rect 2317 25171 2375 25177
rect 6362 25168 6368 25220
rect 6420 25217 6426 25220
rect 6420 25211 6483 25217
rect 6420 25177 6437 25211
rect 6471 25177 6483 25211
rect 6420 25171 6483 25177
rect 6641 25211 6699 25217
rect 6641 25177 6653 25211
rect 6687 25208 6699 25211
rect 6822 25208 6828 25220
rect 6687 25180 6828 25208
rect 6687 25177 6699 25180
rect 6641 25171 6699 25177
rect 6420 25168 6426 25171
rect 6822 25168 6828 25180
rect 6880 25168 6886 25220
rect 8294 25168 8300 25220
rect 8352 25168 8358 25220
rect 1946 25100 1952 25152
rect 2004 25100 2010 25152
rect 2133 25143 2191 25149
rect 2133 25109 2145 25143
rect 2179 25140 2191 25143
rect 2222 25140 2228 25152
rect 2179 25112 2228 25140
rect 2179 25109 2191 25112
rect 2133 25103 2191 25109
rect 2222 25100 2228 25112
rect 2280 25100 2286 25152
rect 5721 25143 5779 25149
rect 5721 25109 5733 25143
rect 5767 25140 5779 25143
rect 6730 25140 6736 25152
rect 5767 25112 6736 25140
rect 5767 25109 5779 25112
rect 5721 25103 5779 25109
rect 6730 25100 6736 25112
rect 6788 25100 6794 25152
rect 8113 25143 8171 25149
rect 8113 25109 8125 25143
rect 8159 25140 8171 25143
rect 8202 25140 8208 25152
rect 8159 25112 8208 25140
rect 8159 25109 8171 25112
rect 8113 25103 8171 25109
rect 8202 25100 8208 25112
rect 8260 25100 8266 25152
rect 1104 25050 19019 25072
rect 1104 24998 5388 25050
rect 5440 24998 5452 25050
rect 5504 24998 5516 25050
rect 5568 24998 5580 25050
rect 5632 24998 5644 25050
rect 5696 24998 9827 25050
rect 9879 24998 9891 25050
rect 9943 24998 9955 25050
rect 10007 24998 10019 25050
rect 10071 24998 10083 25050
rect 10135 24998 14266 25050
rect 14318 24998 14330 25050
rect 14382 24998 14394 25050
rect 14446 24998 14458 25050
rect 14510 24998 14522 25050
rect 14574 24998 18705 25050
rect 18757 24998 18769 25050
rect 18821 24998 18833 25050
rect 18885 24998 18897 25050
rect 18949 24998 18961 25050
rect 19013 24998 19019 25050
rect 1104 24976 19019 24998
rect 3881 24939 3939 24945
rect 3881 24905 3893 24939
rect 3927 24936 3939 24939
rect 4062 24936 4068 24948
rect 3927 24908 4068 24936
rect 3927 24905 3939 24908
rect 3881 24899 3939 24905
rect 4062 24896 4068 24908
rect 4120 24896 4126 24948
rect 5074 24896 5080 24948
rect 5132 24936 5138 24948
rect 5261 24939 5319 24945
rect 5261 24936 5273 24939
rect 5132 24908 5273 24936
rect 5132 24896 5138 24908
rect 5261 24905 5273 24908
rect 5307 24905 5319 24939
rect 5261 24899 5319 24905
rect 6822 24828 6828 24880
rect 6880 24868 6886 24880
rect 7913 24871 7971 24877
rect 6880 24840 7052 24868
rect 6880 24828 6886 24840
rect 4890 24760 4896 24812
rect 4948 24800 4954 24812
rect 7024 24809 7052 24840
rect 7913 24837 7925 24871
rect 7959 24868 7971 24871
rect 8113 24871 8171 24877
rect 7959 24837 7972 24868
rect 7913 24831 7972 24837
rect 8113 24837 8125 24871
rect 8159 24868 8171 24871
rect 8386 24868 8392 24880
rect 8159 24840 8392 24868
rect 8159 24837 8171 24840
rect 8113 24831 8171 24837
rect 5169 24803 5227 24809
rect 5169 24800 5181 24803
rect 4948 24772 5181 24800
rect 4948 24760 4954 24772
rect 5169 24769 5181 24772
rect 5215 24769 5227 24803
rect 5169 24763 5227 24769
rect 5445 24803 5503 24809
rect 5445 24769 5457 24803
rect 5491 24800 5503 24803
rect 6733 24803 6791 24809
rect 5491 24772 6592 24800
rect 5491 24769 5503 24772
rect 5445 24763 5503 24769
rect 2222 24692 2228 24744
rect 2280 24732 2286 24744
rect 3513 24735 3571 24741
rect 3513 24732 3525 24735
rect 2280 24704 3525 24732
rect 2280 24692 2286 24704
rect 3513 24701 3525 24704
rect 3559 24732 3571 24735
rect 4798 24732 4804 24744
rect 3559 24704 4804 24732
rect 3559 24701 3571 24704
rect 3513 24695 3571 24701
rect 4798 24692 4804 24704
rect 4856 24692 4862 24744
rect 6564 24673 6592 24772
rect 6733 24769 6745 24803
rect 6779 24800 6791 24803
rect 7009 24803 7067 24809
rect 6779 24772 6960 24800
rect 6779 24769 6791 24772
rect 6733 24763 6791 24769
rect 6638 24692 6644 24744
rect 6696 24732 6702 24744
rect 6825 24735 6883 24741
rect 6825 24732 6837 24735
rect 6696 24704 6837 24732
rect 6696 24692 6702 24704
rect 6825 24701 6837 24704
rect 6871 24701 6883 24735
rect 6932 24732 6960 24772
rect 7009 24769 7021 24803
rect 7055 24769 7067 24803
rect 7944 24800 7972 24831
rect 8386 24828 8392 24840
rect 8444 24868 8450 24880
rect 9122 24868 9128 24880
rect 8444 24840 9128 24868
rect 8444 24828 8450 24840
rect 9122 24828 9128 24840
rect 9180 24828 9186 24880
rect 8018 24800 8024 24812
rect 7944 24772 8024 24800
rect 7009 24763 7067 24769
rect 8018 24760 8024 24772
rect 8076 24760 8082 24812
rect 7926 24732 7932 24744
rect 6932 24704 7932 24732
rect 6825 24695 6883 24701
rect 7926 24692 7932 24704
rect 7984 24692 7990 24744
rect 4065 24667 4123 24673
rect 4065 24664 4077 24667
rect 3620 24636 4077 24664
rect 2682 24556 2688 24608
rect 2740 24596 2746 24608
rect 3620 24596 3648 24636
rect 4065 24633 4077 24636
rect 4111 24633 4123 24667
rect 4065 24627 4123 24633
rect 6549 24667 6607 24673
rect 6549 24633 6561 24667
rect 6595 24633 6607 24667
rect 6549 24627 6607 24633
rect 7098 24624 7104 24676
rect 7156 24664 7162 24676
rect 7745 24667 7803 24673
rect 7745 24664 7757 24667
rect 7156 24636 7757 24664
rect 7156 24624 7162 24636
rect 7745 24633 7757 24636
rect 7791 24633 7803 24667
rect 7745 24627 7803 24633
rect 2740 24568 3648 24596
rect 3881 24599 3939 24605
rect 2740 24556 2746 24568
rect 3881 24565 3893 24599
rect 3927 24596 3939 24599
rect 4154 24596 4160 24608
rect 3927 24568 4160 24596
rect 3927 24565 3939 24568
rect 3881 24559 3939 24565
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 7009 24599 7067 24605
rect 7009 24565 7021 24599
rect 7055 24596 7067 24599
rect 7466 24596 7472 24608
rect 7055 24568 7472 24596
rect 7055 24565 7067 24568
rect 7009 24559 7067 24565
rect 7466 24556 7472 24568
rect 7524 24556 7530 24608
rect 7558 24556 7564 24608
rect 7616 24596 7622 24608
rect 7929 24599 7987 24605
rect 7929 24596 7941 24599
rect 7616 24568 7941 24596
rect 7616 24556 7622 24568
rect 7929 24565 7941 24568
rect 7975 24565 7987 24599
rect 7929 24559 7987 24565
rect 1104 24506 18860 24528
rect 1104 24454 3169 24506
rect 3221 24454 3233 24506
rect 3285 24454 3297 24506
rect 3349 24454 3361 24506
rect 3413 24454 3425 24506
rect 3477 24454 7608 24506
rect 7660 24454 7672 24506
rect 7724 24454 7736 24506
rect 7788 24454 7800 24506
rect 7852 24454 7864 24506
rect 7916 24454 12047 24506
rect 12099 24454 12111 24506
rect 12163 24454 12175 24506
rect 12227 24454 12239 24506
rect 12291 24454 12303 24506
rect 12355 24454 16486 24506
rect 16538 24454 16550 24506
rect 16602 24454 16614 24506
rect 16666 24454 16678 24506
rect 16730 24454 16742 24506
rect 16794 24454 18860 24506
rect 1104 24432 18860 24454
rect 4154 24352 4160 24404
rect 4212 24352 4218 24404
rect 5629 24395 5687 24401
rect 5629 24392 5641 24395
rect 4264 24364 5641 24392
rect 2222 24256 2228 24268
rect 1872 24228 2228 24256
rect 1872 24197 1900 24228
rect 2222 24216 2228 24228
rect 2280 24216 2286 24268
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24157 1915 24191
rect 1857 24151 1915 24157
rect 2130 24148 2136 24200
rect 2188 24148 2194 24200
rect 4264 24188 4292 24364
rect 5629 24361 5641 24364
rect 5675 24392 5687 24395
rect 6270 24392 6276 24404
rect 5675 24364 6276 24392
rect 5675 24361 5687 24364
rect 5629 24355 5687 24361
rect 6270 24352 6276 24364
rect 6328 24392 6334 24404
rect 6730 24392 6736 24404
rect 6328 24364 6736 24392
rect 6328 24352 6334 24364
rect 6730 24352 6736 24364
rect 6788 24392 6794 24404
rect 7834 24392 7840 24404
rect 6788 24364 7840 24392
rect 6788 24352 6794 24364
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 5810 24324 5816 24336
rect 4356 24296 5816 24324
rect 4356 24265 4384 24296
rect 5810 24284 5816 24296
rect 5868 24324 5874 24336
rect 8021 24327 8079 24333
rect 8021 24324 8033 24327
rect 5868 24296 8033 24324
rect 5868 24284 5874 24296
rect 4341 24259 4399 24265
rect 4341 24225 4353 24259
rect 4387 24225 4399 24259
rect 4341 24219 4399 24225
rect 4525 24259 4583 24265
rect 4525 24225 4537 24259
rect 4571 24256 4583 24259
rect 4571 24228 5028 24256
rect 4571 24225 4583 24228
rect 4525 24219 4583 24225
rect 5000 24200 5028 24228
rect 4433 24191 4491 24197
rect 4433 24188 4445 24191
rect 4264 24160 4445 24188
rect 4433 24157 4445 24160
rect 4479 24157 4491 24191
rect 4433 24151 4491 24157
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 1026 24080 1032 24132
rect 1084 24120 1090 24132
rect 2148 24120 2176 24148
rect 1084 24092 2176 24120
rect 4632 24120 4660 24151
rect 4982 24148 4988 24200
rect 5040 24188 5046 24200
rect 5169 24191 5227 24197
rect 5169 24188 5181 24191
rect 5040 24160 5181 24188
rect 5040 24148 5046 24160
rect 5169 24157 5181 24160
rect 5215 24157 5227 24191
rect 5169 24151 5227 24157
rect 5537 24191 5595 24197
rect 5537 24157 5549 24191
rect 5583 24157 5595 24191
rect 5537 24151 5595 24157
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24188 5779 24191
rect 6012 24188 6040 24296
rect 8021 24293 8033 24296
rect 8067 24293 8079 24327
rect 8021 24287 8079 24293
rect 7006 24216 7012 24268
rect 7064 24256 7070 24268
rect 7064 24228 8248 24256
rect 7064 24216 7070 24228
rect 6086 24188 6092 24200
rect 5767 24160 6092 24188
rect 5767 24157 5779 24160
rect 5721 24151 5779 24157
rect 5552 24120 5580 24151
rect 6086 24148 6092 24160
rect 6144 24148 6150 24200
rect 6546 24148 6552 24200
rect 6604 24188 6610 24200
rect 6917 24191 6975 24197
rect 6917 24188 6929 24191
rect 6604 24160 6929 24188
rect 6604 24148 6610 24160
rect 6917 24157 6929 24160
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 7282 24148 7288 24200
rect 7340 24188 7346 24200
rect 7377 24191 7435 24197
rect 7377 24188 7389 24191
rect 7340 24160 7389 24188
rect 7340 24148 7346 24160
rect 7377 24157 7389 24160
rect 7423 24157 7435 24191
rect 7377 24151 7435 24157
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 8220 24197 8248 24228
rect 7929 24191 7987 24197
rect 7929 24188 7941 24191
rect 7892 24160 7941 24188
rect 7892 24148 7898 24160
rect 7929 24157 7941 24160
rect 7975 24157 7987 24191
rect 7929 24151 7987 24157
rect 8205 24191 8263 24197
rect 8205 24157 8217 24191
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 5810 24120 5816 24132
rect 4632 24092 5816 24120
rect 1084 24080 1090 24092
rect 5810 24080 5816 24092
rect 5868 24080 5874 24132
rect 7193 24123 7251 24129
rect 7193 24089 7205 24123
rect 7239 24120 7251 24123
rect 9674 24120 9680 24132
rect 7239 24092 9680 24120
rect 7239 24089 7251 24092
rect 7193 24083 7251 24089
rect 9674 24080 9680 24092
rect 9732 24080 9738 24132
rect 1949 24055 2007 24061
rect 1949 24021 1961 24055
rect 1995 24052 2007 24055
rect 2038 24052 2044 24064
rect 1995 24024 2044 24052
rect 1995 24021 2007 24024
rect 1949 24015 2007 24021
rect 2038 24012 2044 24024
rect 2096 24012 2102 24064
rect 2317 24055 2375 24061
rect 2317 24021 2329 24055
rect 2363 24052 2375 24055
rect 2958 24052 2964 24064
rect 2363 24024 2964 24052
rect 2363 24021 2375 24024
rect 2317 24015 2375 24021
rect 2958 24012 2964 24024
rect 3016 24012 3022 24064
rect 4338 24012 4344 24064
rect 4396 24052 4402 24064
rect 5353 24055 5411 24061
rect 5353 24052 5365 24055
rect 4396 24024 5365 24052
rect 4396 24012 4402 24024
rect 5353 24021 5365 24024
rect 5399 24021 5411 24055
rect 5353 24015 5411 24021
rect 8389 24055 8447 24061
rect 8389 24021 8401 24055
rect 8435 24052 8447 24055
rect 9030 24052 9036 24064
rect 8435 24024 9036 24052
rect 8435 24021 8447 24024
rect 8389 24015 8447 24021
rect 9030 24012 9036 24024
rect 9088 24012 9094 24064
rect 1104 23962 19019 23984
rect 1104 23910 5388 23962
rect 5440 23910 5452 23962
rect 5504 23910 5516 23962
rect 5568 23910 5580 23962
rect 5632 23910 5644 23962
rect 5696 23910 9827 23962
rect 9879 23910 9891 23962
rect 9943 23910 9955 23962
rect 10007 23910 10019 23962
rect 10071 23910 10083 23962
rect 10135 23910 14266 23962
rect 14318 23910 14330 23962
rect 14382 23910 14394 23962
rect 14446 23910 14458 23962
rect 14510 23910 14522 23962
rect 14574 23910 18705 23962
rect 18757 23910 18769 23962
rect 18821 23910 18833 23962
rect 18885 23910 18897 23962
rect 18949 23910 18961 23962
rect 19013 23910 19019 23962
rect 1104 23888 19019 23910
rect 4062 23808 4068 23860
rect 4120 23808 4126 23860
rect 4338 23808 4344 23860
rect 4396 23848 4402 23860
rect 4706 23848 4712 23860
rect 4396 23820 4712 23848
rect 4396 23808 4402 23820
rect 4706 23808 4712 23820
rect 4764 23808 4770 23860
rect 6362 23808 6368 23860
rect 6420 23848 6426 23860
rect 7561 23851 7619 23857
rect 7561 23848 7573 23851
rect 6420 23820 7573 23848
rect 6420 23808 6426 23820
rect 7561 23817 7573 23820
rect 7607 23817 7619 23851
rect 7561 23811 7619 23817
rect 4080 23780 4108 23808
rect 4080 23752 7144 23780
rect 7116 23724 7144 23752
rect 4062 23672 4068 23724
rect 4120 23672 4126 23724
rect 4246 23672 4252 23724
rect 4304 23672 4310 23724
rect 4706 23672 4712 23724
rect 4764 23712 4770 23724
rect 5258 23712 5264 23724
rect 4764 23684 5264 23712
rect 4764 23672 4770 23684
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 7098 23672 7104 23724
rect 7156 23672 7162 23724
rect 7466 23672 7472 23724
rect 7524 23712 7530 23724
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 7524 23684 7757 23712
rect 7524 23672 7530 23684
rect 7745 23681 7757 23684
rect 7791 23681 7803 23715
rect 7745 23675 7803 23681
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 6546 23604 6552 23656
rect 6604 23644 6610 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6604 23616 6837 23644
rect 6604 23604 6610 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 6825 23607 6883 23613
rect 4246 23536 4252 23588
rect 4304 23576 4310 23588
rect 4341 23579 4399 23585
rect 4341 23576 4353 23579
rect 4304 23548 4353 23576
rect 4304 23536 4310 23548
rect 4341 23545 4353 23548
rect 4387 23545 4399 23579
rect 4341 23539 4399 23545
rect 934 23468 940 23520
rect 992 23508 998 23520
rect 1581 23511 1639 23517
rect 1581 23508 1593 23511
rect 992 23480 1593 23508
rect 992 23468 998 23480
rect 1581 23477 1593 23480
rect 1627 23477 1639 23511
rect 1581 23471 1639 23477
rect 1104 23418 18860 23440
rect 1104 23366 3169 23418
rect 3221 23366 3233 23418
rect 3285 23366 3297 23418
rect 3349 23366 3361 23418
rect 3413 23366 3425 23418
rect 3477 23366 7608 23418
rect 7660 23366 7672 23418
rect 7724 23366 7736 23418
rect 7788 23366 7800 23418
rect 7852 23366 7864 23418
rect 7916 23366 12047 23418
rect 12099 23366 12111 23418
rect 12163 23366 12175 23418
rect 12227 23366 12239 23418
rect 12291 23366 12303 23418
rect 12355 23366 16486 23418
rect 16538 23366 16550 23418
rect 16602 23366 16614 23418
rect 16666 23366 16678 23418
rect 16730 23366 16742 23418
rect 16794 23366 18860 23418
rect 1104 23344 18860 23366
rect 5902 23264 5908 23316
rect 5960 23264 5966 23316
rect 6825 23307 6883 23313
rect 6825 23273 6837 23307
rect 6871 23304 6883 23307
rect 8294 23304 8300 23316
rect 6871 23276 8300 23304
rect 6871 23273 6883 23276
rect 6825 23267 6883 23273
rect 5813 23239 5871 23245
rect 5813 23205 5825 23239
rect 5859 23236 5871 23239
rect 5994 23236 6000 23248
rect 5859 23208 6000 23236
rect 5859 23205 5871 23208
rect 5813 23199 5871 23205
rect 5994 23196 6000 23208
rect 6052 23196 6058 23248
rect 5721 23171 5779 23177
rect 5721 23137 5733 23171
rect 5767 23168 5779 23171
rect 6178 23168 6184 23180
rect 5767 23140 6184 23168
rect 5767 23137 5779 23140
rect 5721 23131 5779 23137
rect 6178 23128 6184 23140
rect 6236 23168 6242 23180
rect 6840 23168 6868 23267
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 6236 23140 6868 23168
rect 6236 23128 6242 23140
rect 5994 23060 6000 23112
rect 6052 23060 6058 23112
rect 6546 22992 6552 23044
rect 6604 22992 6610 23044
rect 7098 22924 7104 22976
rect 7156 22964 7162 22976
rect 8294 22964 8300 22976
rect 7156 22936 8300 22964
rect 7156 22924 7162 22936
rect 8294 22924 8300 22936
rect 8352 22924 8358 22976
rect 1104 22874 19019 22896
rect 1104 22822 5388 22874
rect 5440 22822 5452 22874
rect 5504 22822 5516 22874
rect 5568 22822 5580 22874
rect 5632 22822 5644 22874
rect 5696 22822 9827 22874
rect 9879 22822 9891 22874
rect 9943 22822 9955 22874
rect 10007 22822 10019 22874
rect 10071 22822 10083 22874
rect 10135 22822 14266 22874
rect 14318 22822 14330 22874
rect 14382 22822 14394 22874
rect 14446 22822 14458 22874
rect 14510 22822 14522 22874
rect 14574 22822 18705 22874
rect 18757 22822 18769 22874
rect 18821 22822 18833 22874
rect 18885 22822 18897 22874
rect 18949 22822 18961 22874
rect 19013 22822 19019 22874
rect 1104 22800 19019 22822
rect 5718 22720 5724 22772
rect 5776 22720 5782 22772
rect 5813 22763 5871 22769
rect 5813 22729 5825 22763
rect 5859 22760 5871 22763
rect 5994 22760 6000 22772
rect 5859 22732 6000 22760
rect 5859 22729 5871 22732
rect 5813 22723 5871 22729
rect 5994 22720 6000 22732
rect 6052 22760 6058 22772
rect 6822 22760 6828 22772
rect 6052 22732 6828 22760
rect 6052 22720 6058 22732
rect 6822 22720 6828 22732
rect 6880 22760 6886 22772
rect 7282 22760 7288 22772
rect 6880 22732 7288 22760
rect 6880 22720 6886 22732
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 7469 22763 7527 22769
rect 7469 22729 7481 22763
rect 7515 22760 7527 22763
rect 8110 22760 8116 22772
rect 7515 22732 8116 22760
rect 7515 22729 7527 22732
rect 7469 22723 7527 22729
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 8205 22763 8263 22769
rect 8205 22729 8217 22763
rect 8251 22760 8263 22763
rect 8294 22760 8300 22772
rect 8251 22732 8300 22760
rect 8251 22729 8263 22732
rect 8205 22723 8263 22729
rect 8294 22720 8300 22732
rect 8352 22720 8358 22772
rect 1762 22692 1768 22704
rect 1596 22664 1768 22692
rect 1596 22633 1624 22664
rect 1762 22652 1768 22664
rect 1820 22692 1826 22704
rect 2590 22692 2596 22704
rect 1820 22664 2596 22692
rect 1820 22652 1826 22664
rect 2590 22652 2596 22664
rect 2648 22652 2654 22704
rect 4062 22652 4068 22704
rect 4120 22692 4126 22704
rect 5261 22695 5319 22701
rect 5261 22692 5273 22695
rect 4120 22664 5273 22692
rect 4120 22652 4126 22664
rect 5261 22661 5273 22664
rect 5307 22661 5319 22695
rect 5261 22655 5319 22661
rect 5629 22695 5687 22701
rect 5629 22661 5641 22695
rect 5675 22692 5687 22695
rect 6362 22692 6368 22704
rect 5675 22664 6368 22692
rect 5675 22661 5687 22664
rect 5629 22655 5687 22661
rect 6362 22652 6368 22664
rect 6420 22652 6426 22704
rect 7374 22652 7380 22704
rect 7432 22692 7438 22704
rect 7432 22664 7972 22692
rect 7432 22652 7438 22664
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22593 1639 22627
rect 1581 22587 1639 22593
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 1946 22624 1952 22636
rect 1719 22596 1952 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 1946 22584 1952 22596
rect 2004 22584 2010 22636
rect 5994 22584 6000 22636
rect 6052 22624 6058 22636
rect 6638 22624 6644 22636
rect 6052 22596 6644 22624
rect 6052 22584 6058 22596
rect 6638 22584 6644 22596
rect 6696 22584 6702 22636
rect 7098 22584 7104 22636
rect 7156 22584 7162 22636
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22624 7343 22627
rect 7466 22624 7472 22636
rect 7331 22596 7472 22624
rect 7331 22593 7343 22596
rect 7285 22587 7343 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 1854 22516 1860 22568
rect 1912 22516 1918 22568
rect 7944 22432 7972 22664
rect 8294 22584 8300 22636
rect 8352 22584 8358 22636
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22624 8539 22627
rect 8938 22624 8944 22636
rect 8527 22596 8944 22624
rect 8527 22593 8539 22596
rect 8481 22587 8539 22593
rect 8938 22584 8944 22596
rect 8996 22584 9002 22636
rect 1765 22423 1823 22429
rect 1765 22389 1777 22423
rect 1811 22420 1823 22423
rect 2130 22420 2136 22432
rect 1811 22392 2136 22420
rect 1811 22389 1823 22392
rect 1765 22383 1823 22389
rect 2130 22380 2136 22392
rect 2188 22380 2194 22432
rect 7466 22380 7472 22432
rect 7524 22420 7530 22432
rect 7834 22420 7840 22432
rect 7524 22392 7840 22420
rect 7524 22380 7530 22392
rect 7834 22380 7840 22392
rect 7892 22380 7898 22432
rect 7926 22380 7932 22432
rect 7984 22380 7990 22432
rect 1104 22330 18860 22352
rect 1104 22278 3169 22330
rect 3221 22278 3233 22330
rect 3285 22278 3297 22330
rect 3349 22278 3361 22330
rect 3413 22278 3425 22330
rect 3477 22278 7608 22330
rect 7660 22278 7672 22330
rect 7724 22278 7736 22330
rect 7788 22278 7800 22330
rect 7852 22278 7864 22330
rect 7916 22278 12047 22330
rect 12099 22278 12111 22330
rect 12163 22278 12175 22330
rect 12227 22278 12239 22330
rect 12291 22278 12303 22330
rect 12355 22278 16486 22330
rect 16538 22278 16550 22330
rect 16602 22278 16614 22330
rect 16666 22278 16678 22330
rect 16730 22278 16742 22330
rect 16794 22278 18860 22330
rect 1104 22256 18860 22278
rect 4430 22176 4436 22228
rect 4488 22176 4494 22228
rect 5718 22176 5724 22228
rect 5776 22216 5782 22228
rect 7098 22216 7104 22228
rect 5776 22188 7104 22216
rect 5776 22176 5782 22188
rect 7098 22176 7104 22188
rect 7156 22176 7162 22228
rect 7190 22176 7196 22228
rect 7248 22216 7254 22228
rect 8110 22216 8116 22228
rect 7248 22188 8116 22216
rect 7248 22176 7254 22188
rect 8110 22176 8116 22188
rect 8168 22176 8174 22228
rect 6178 22080 6184 22092
rect 4632 22052 6184 22080
rect 1854 21904 1860 21956
rect 1912 21944 1918 21956
rect 2774 21944 2780 21956
rect 1912 21916 2780 21944
rect 1912 21904 1918 21916
rect 2774 21904 2780 21916
rect 2832 21944 2838 21956
rect 4632 21953 4660 22052
rect 6178 22040 6184 22052
rect 6236 22040 6242 22092
rect 4982 21972 4988 22024
rect 5040 22012 5046 22024
rect 5629 22015 5687 22021
rect 5629 22012 5641 22015
rect 5040 21984 5641 22012
rect 5040 21972 5046 21984
rect 5629 21981 5641 21984
rect 5675 21981 5687 22015
rect 6086 22012 6092 22024
rect 5629 21975 5687 21981
rect 5736 21984 6092 22012
rect 5736 21956 5764 21984
rect 6086 21972 6092 21984
rect 6144 21972 6150 22024
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 7156 21984 7481 22012
rect 7156 21972 7162 21984
rect 7469 21981 7481 21984
rect 7515 21981 7527 22015
rect 7469 21975 7527 21981
rect 7653 22015 7711 22021
rect 7653 21981 7665 22015
rect 7699 21981 7711 22015
rect 7653 21975 7711 21981
rect 4617 21947 4675 21953
rect 4617 21944 4629 21947
rect 2832 21916 4629 21944
rect 2832 21904 2838 21916
rect 4617 21913 4629 21916
rect 4663 21913 4675 21947
rect 4617 21907 4675 21913
rect 4798 21904 4804 21956
rect 4856 21944 4862 21956
rect 5077 21947 5135 21953
rect 5077 21944 5089 21947
rect 4856 21916 5089 21944
rect 4856 21904 4862 21916
rect 5077 21913 5089 21916
rect 5123 21913 5135 21947
rect 5077 21907 5135 21913
rect 5445 21947 5503 21953
rect 5445 21913 5457 21947
rect 5491 21944 5503 21947
rect 5718 21944 5724 21956
rect 5491 21916 5724 21944
rect 5491 21913 5503 21916
rect 5445 21907 5503 21913
rect 5718 21904 5724 21916
rect 5776 21904 5782 21956
rect 5810 21904 5816 21956
rect 5868 21944 5874 21956
rect 6178 21944 6184 21956
rect 5868 21916 6184 21944
rect 5868 21904 5874 21916
rect 6178 21904 6184 21916
rect 6236 21904 6242 21956
rect 7374 21904 7380 21956
rect 7432 21944 7438 21956
rect 7668 21944 7696 21975
rect 7432 21916 7696 21944
rect 7432 21904 7438 21916
rect 7834 21904 7840 21956
rect 7892 21944 7898 21956
rect 8202 21944 8208 21956
rect 7892 21916 8208 21944
rect 7892 21904 7898 21916
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 1578 21836 1584 21888
rect 1636 21876 1642 21888
rect 4249 21879 4307 21885
rect 4249 21876 4261 21879
rect 1636 21848 4261 21876
rect 1636 21836 1642 21848
rect 4249 21845 4261 21848
rect 4295 21845 4307 21879
rect 4249 21839 4307 21845
rect 4417 21879 4475 21885
rect 4417 21845 4429 21879
rect 4463 21876 4475 21879
rect 5258 21876 5264 21888
rect 4463 21848 5264 21876
rect 4463 21845 4475 21848
rect 4417 21839 4475 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 5537 21879 5595 21885
rect 5537 21845 5549 21879
rect 5583 21876 5595 21879
rect 6086 21876 6092 21888
rect 5583 21848 6092 21876
rect 5583 21845 5595 21848
rect 5537 21839 5595 21845
rect 6086 21836 6092 21848
rect 6144 21876 6150 21888
rect 6362 21876 6368 21888
rect 6144 21848 6368 21876
rect 6144 21836 6150 21848
rect 6362 21836 6368 21848
rect 6420 21836 6426 21888
rect 1104 21786 19019 21808
rect 1104 21734 5388 21786
rect 5440 21734 5452 21786
rect 5504 21734 5516 21786
rect 5568 21734 5580 21786
rect 5632 21734 5644 21786
rect 5696 21734 9827 21786
rect 9879 21734 9891 21786
rect 9943 21734 9955 21786
rect 10007 21734 10019 21786
rect 10071 21734 10083 21786
rect 10135 21734 14266 21786
rect 14318 21734 14330 21786
rect 14382 21734 14394 21786
rect 14446 21734 14458 21786
rect 14510 21734 14522 21786
rect 14574 21734 18705 21786
rect 18757 21734 18769 21786
rect 18821 21734 18833 21786
rect 18885 21734 18897 21786
rect 18949 21734 18961 21786
rect 19013 21734 19019 21786
rect 1104 21712 19019 21734
rect 5258 21632 5264 21684
rect 5316 21672 5322 21684
rect 5353 21675 5411 21681
rect 5353 21672 5365 21675
rect 5316 21644 5365 21672
rect 5316 21632 5322 21644
rect 5353 21641 5365 21644
rect 5399 21641 5411 21675
rect 6086 21672 6092 21684
rect 5353 21635 5411 21641
rect 5736 21644 6092 21672
rect 5736 21548 5764 21644
rect 6086 21632 6092 21644
rect 6144 21632 6150 21684
rect 5902 21564 5908 21616
rect 5960 21604 5966 21616
rect 5960 21576 7788 21604
rect 5960 21564 5966 21576
rect 4982 21496 4988 21548
rect 5040 21536 5046 21548
rect 5258 21536 5264 21548
rect 5040 21508 5264 21536
rect 5040 21496 5046 21508
rect 5258 21496 5264 21508
rect 5316 21536 5322 21548
rect 5537 21539 5595 21545
rect 5537 21536 5549 21539
rect 5316 21508 5549 21536
rect 5316 21496 5322 21508
rect 5537 21505 5549 21508
rect 5583 21505 5595 21539
rect 5537 21499 5595 21505
rect 5718 21496 5724 21548
rect 5776 21496 5782 21548
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 7285 21539 7343 21545
rect 7285 21505 7297 21539
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7760 21536 7788 21576
rect 7834 21564 7840 21616
rect 7892 21604 7898 21616
rect 7892 21576 8800 21604
rect 7892 21564 7898 21576
rect 8021 21539 8079 21545
rect 8021 21536 8033 21539
rect 7760 21508 8033 21536
rect 7653 21499 7711 21505
rect 8021 21505 8033 21508
rect 8067 21505 8079 21539
rect 8021 21499 8079 21505
rect 5902 21428 5908 21480
rect 5960 21468 5966 21480
rect 7300 21468 7328 21499
rect 5960 21440 7328 21468
rect 7668 21468 7696 21499
rect 8202 21496 8208 21548
rect 8260 21536 8266 21548
rect 8772 21545 8800 21576
rect 8389 21539 8447 21545
rect 8389 21536 8401 21539
rect 8260 21508 8401 21536
rect 8260 21496 8266 21508
rect 8389 21505 8401 21508
rect 8435 21505 8447 21539
rect 8389 21499 8447 21505
rect 8757 21539 8815 21545
rect 8757 21505 8769 21539
rect 8803 21505 8815 21539
rect 8757 21499 8815 21505
rect 8938 21468 8944 21480
rect 7668 21440 8944 21468
rect 5960 21428 5966 21440
rect 7300 21332 7328 21440
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 7469 21403 7527 21409
rect 7469 21369 7481 21403
rect 7515 21400 7527 21403
rect 8386 21400 8392 21412
rect 7515 21372 8392 21400
rect 7515 21369 7527 21372
rect 7469 21363 7527 21369
rect 8386 21360 8392 21372
rect 8444 21360 8450 21412
rect 8294 21332 8300 21344
rect 7300 21304 8300 21332
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 1104 21242 18860 21264
rect 1104 21190 3169 21242
rect 3221 21190 3233 21242
rect 3285 21190 3297 21242
rect 3349 21190 3361 21242
rect 3413 21190 3425 21242
rect 3477 21190 7608 21242
rect 7660 21190 7672 21242
rect 7724 21190 7736 21242
rect 7788 21190 7800 21242
rect 7852 21190 7864 21242
rect 7916 21190 12047 21242
rect 12099 21190 12111 21242
rect 12163 21190 12175 21242
rect 12227 21190 12239 21242
rect 12291 21190 12303 21242
rect 12355 21190 16486 21242
rect 16538 21190 16550 21242
rect 16602 21190 16614 21242
rect 16666 21190 16678 21242
rect 16730 21190 16742 21242
rect 16794 21190 18860 21242
rect 1104 21168 18860 21190
rect 2041 21131 2099 21137
rect 2041 21097 2053 21131
rect 2087 21128 2099 21131
rect 2222 21128 2228 21140
rect 2087 21100 2228 21128
rect 2087 21097 2099 21100
rect 2041 21091 2099 21097
rect 2222 21088 2228 21100
rect 2280 21088 2286 21140
rect 5074 21088 5080 21140
rect 5132 21088 5138 21140
rect 8202 21088 8208 21140
rect 8260 21088 8266 21140
rect 1857 20995 1915 21001
rect 1857 20961 1869 20995
rect 1903 20992 1915 20995
rect 2774 20992 2780 21004
rect 1903 20964 2780 20992
rect 1903 20961 1915 20964
rect 1857 20955 1915 20961
rect 2774 20952 2780 20964
rect 2832 20992 2838 21004
rect 2869 20995 2927 21001
rect 2869 20992 2881 20995
rect 2832 20964 2881 20992
rect 2832 20952 2838 20964
rect 2869 20961 2881 20964
rect 2915 20961 2927 20995
rect 2869 20955 2927 20961
rect 2038 20884 2044 20936
rect 2096 20924 2102 20936
rect 2133 20927 2191 20933
rect 2133 20924 2145 20927
rect 2096 20896 2145 20924
rect 2096 20884 2102 20896
rect 2133 20893 2145 20896
rect 2179 20924 2191 20927
rect 2222 20924 2228 20936
rect 2179 20896 2228 20924
rect 2179 20893 2191 20896
rect 2133 20887 2191 20893
rect 2222 20884 2228 20896
rect 2280 20884 2286 20936
rect 3329 20927 3387 20933
rect 3329 20893 3341 20927
rect 3375 20924 3387 20927
rect 3694 20924 3700 20936
rect 3375 20896 3700 20924
rect 3375 20893 3387 20896
rect 3329 20887 3387 20893
rect 3694 20884 3700 20896
rect 3752 20884 3758 20936
rect 5166 20884 5172 20936
rect 5224 20924 5230 20936
rect 5353 20927 5411 20933
rect 5353 20924 5365 20927
rect 5224 20896 5365 20924
rect 5224 20884 5230 20896
rect 5353 20893 5365 20896
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 7466 20884 7472 20936
rect 7524 20924 7530 20936
rect 8113 20927 8171 20933
rect 8113 20924 8125 20927
rect 7524 20896 8125 20924
rect 7524 20884 7530 20896
rect 8113 20893 8125 20896
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 3050 20816 3056 20868
rect 3108 20856 3114 20868
rect 3237 20859 3295 20865
rect 3237 20856 3249 20859
rect 3108 20828 3249 20856
rect 3108 20816 3114 20828
rect 3237 20825 3249 20828
rect 3283 20825 3295 20859
rect 3237 20819 3295 20825
rect 3970 20816 3976 20868
rect 4028 20856 4034 20868
rect 5261 20859 5319 20865
rect 5261 20856 5273 20859
rect 4028 20828 5273 20856
rect 4028 20816 4034 20828
rect 5261 20825 5273 20828
rect 5307 20825 5319 20859
rect 5261 20819 5319 20825
rect 5813 20859 5871 20865
rect 5813 20825 5825 20859
rect 5859 20856 5871 20859
rect 5902 20856 5908 20868
rect 5859 20828 5908 20856
rect 5859 20825 5871 20828
rect 5813 20819 5871 20825
rect 5902 20816 5908 20828
rect 5960 20816 5966 20868
rect 1854 20748 1860 20800
rect 1912 20748 1918 20800
rect 3142 20748 3148 20800
rect 3200 20748 3206 20800
rect 7190 20748 7196 20800
rect 7248 20788 7254 20800
rect 7466 20788 7472 20800
rect 7248 20760 7472 20788
rect 7248 20748 7254 20760
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 1104 20698 19019 20720
rect 1104 20646 5388 20698
rect 5440 20646 5452 20698
rect 5504 20646 5516 20698
rect 5568 20646 5580 20698
rect 5632 20646 5644 20698
rect 5696 20646 9827 20698
rect 9879 20646 9891 20698
rect 9943 20646 9955 20698
rect 10007 20646 10019 20698
rect 10071 20646 10083 20698
rect 10135 20646 14266 20698
rect 14318 20646 14330 20698
rect 14382 20646 14394 20698
rect 14446 20646 14458 20698
rect 14510 20646 14522 20698
rect 14574 20646 18705 20698
rect 18757 20646 18769 20698
rect 18821 20646 18833 20698
rect 18885 20646 18897 20698
rect 18949 20646 18961 20698
rect 19013 20646 19019 20698
rect 1104 20624 19019 20646
rect 4430 20544 4436 20596
rect 4488 20584 4494 20596
rect 5261 20587 5319 20593
rect 5261 20584 5273 20587
rect 4488 20556 5273 20584
rect 4488 20544 4494 20556
rect 5261 20553 5273 20556
rect 5307 20553 5319 20587
rect 5261 20547 5319 20553
rect 5353 20519 5411 20525
rect 5353 20485 5365 20519
rect 5399 20516 5411 20519
rect 5718 20516 5724 20528
rect 5399 20488 5724 20516
rect 5399 20485 5411 20488
rect 5353 20479 5411 20485
rect 5718 20476 5724 20488
rect 5776 20516 5782 20528
rect 6086 20516 6092 20528
rect 5776 20488 6092 20516
rect 5776 20476 5782 20488
rect 6086 20476 6092 20488
rect 6144 20476 6150 20528
rect 3142 20408 3148 20460
rect 3200 20448 3206 20460
rect 3697 20451 3755 20457
rect 3697 20448 3709 20451
rect 3200 20420 3709 20448
rect 3200 20408 3206 20420
rect 3697 20417 3709 20420
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 5258 20408 5264 20460
rect 5316 20408 5322 20460
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20448 5595 20451
rect 5810 20448 5816 20460
rect 5583 20420 5816 20448
rect 5583 20417 5595 20420
rect 5537 20411 5595 20417
rect 5810 20408 5816 20420
rect 5868 20448 5874 20460
rect 6362 20448 6368 20460
rect 5868 20420 6368 20448
rect 5868 20408 5874 20420
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 3050 20340 3056 20392
rect 3108 20380 3114 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3108 20352 3433 20380
rect 3108 20340 3114 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 6270 20340 6276 20392
rect 6328 20380 6334 20392
rect 6546 20380 6552 20392
rect 6328 20352 6552 20380
rect 6328 20340 6334 20352
rect 6546 20340 6552 20352
rect 6604 20340 6610 20392
rect 3513 20247 3571 20253
rect 3513 20213 3525 20247
rect 3559 20244 3571 20247
rect 3694 20244 3700 20256
rect 3559 20216 3700 20244
rect 3559 20213 3571 20216
rect 3513 20207 3571 20213
rect 3694 20204 3700 20216
rect 3752 20204 3758 20256
rect 3881 20247 3939 20253
rect 3881 20213 3893 20247
rect 3927 20244 3939 20247
rect 6546 20244 6552 20256
rect 3927 20216 6552 20244
rect 3927 20213 3939 20216
rect 3881 20207 3939 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 1104 20154 18860 20176
rect 1104 20102 3169 20154
rect 3221 20102 3233 20154
rect 3285 20102 3297 20154
rect 3349 20102 3361 20154
rect 3413 20102 3425 20154
rect 3477 20102 7608 20154
rect 7660 20102 7672 20154
rect 7724 20102 7736 20154
rect 7788 20102 7800 20154
rect 7852 20102 7864 20154
rect 7916 20102 12047 20154
rect 12099 20102 12111 20154
rect 12163 20102 12175 20154
rect 12227 20102 12239 20154
rect 12291 20102 12303 20154
rect 12355 20102 16486 20154
rect 16538 20102 16550 20154
rect 16602 20102 16614 20154
rect 16666 20102 16678 20154
rect 16730 20102 16742 20154
rect 16794 20102 18860 20154
rect 1104 20080 18860 20102
rect 2958 20000 2964 20052
rect 3016 20000 3022 20052
rect 1946 19932 1952 19984
rect 2004 19972 2010 19984
rect 2593 19975 2651 19981
rect 2593 19972 2605 19975
rect 2004 19944 2605 19972
rect 2004 19932 2010 19944
rect 2593 19941 2605 19944
rect 2639 19941 2651 19975
rect 2593 19935 2651 19941
rect 1210 19796 1216 19848
rect 1268 19836 1274 19848
rect 1765 19839 1823 19845
rect 1765 19836 1777 19839
rect 1268 19808 1777 19836
rect 1268 19796 1274 19808
rect 1765 19805 1777 19808
rect 1811 19805 1823 19839
rect 1765 19799 1823 19805
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 1581 19771 1639 19777
rect 1581 19768 1593 19771
rect 992 19740 1593 19768
rect 992 19728 998 19740
rect 1581 19737 1593 19740
rect 1627 19737 1639 19771
rect 1581 19731 1639 19737
rect 2774 19728 2780 19780
rect 2832 19768 2838 19780
rect 2961 19771 3019 19777
rect 2961 19768 2973 19771
rect 2832 19740 2973 19768
rect 2832 19728 2838 19740
rect 2961 19737 2973 19740
rect 3007 19768 3019 19771
rect 3970 19768 3976 19780
rect 3007 19740 3976 19768
rect 3007 19737 3019 19740
rect 2961 19731 3019 19737
rect 3970 19728 3976 19740
rect 4028 19728 4034 19780
rect 3145 19703 3203 19709
rect 3145 19669 3157 19703
rect 3191 19700 3203 19703
rect 4062 19700 4068 19712
rect 3191 19672 4068 19700
rect 3191 19669 3203 19672
rect 3145 19663 3203 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 1104 19610 19019 19632
rect 1104 19558 5388 19610
rect 5440 19558 5452 19610
rect 5504 19558 5516 19610
rect 5568 19558 5580 19610
rect 5632 19558 5644 19610
rect 5696 19558 9827 19610
rect 9879 19558 9891 19610
rect 9943 19558 9955 19610
rect 10007 19558 10019 19610
rect 10071 19558 10083 19610
rect 10135 19558 14266 19610
rect 14318 19558 14330 19610
rect 14382 19558 14394 19610
rect 14446 19558 14458 19610
rect 14510 19558 14522 19610
rect 14574 19558 18705 19610
rect 18757 19558 18769 19610
rect 18821 19558 18833 19610
rect 18885 19558 18897 19610
rect 18949 19558 18961 19610
rect 19013 19558 19019 19610
rect 1104 19536 19019 19558
rect 2783 19499 2841 19505
rect 2783 19465 2795 19499
rect 2829 19496 2841 19499
rect 4430 19496 4436 19508
rect 2829 19468 4436 19496
rect 2829 19465 2841 19468
rect 2783 19459 2841 19465
rect 4430 19456 4436 19468
rect 4488 19456 4494 19508
rect 1854 19388 1860 19440
rect 1912 19428 1918 19440
rect 2685 19431 2743 19437
rect 2685 19428 2697 19431
rect 1912 19400 2697 19428
rect 1912 19388 1918 19400
rect 2685 19397 2697 19400
rect 2731 19397 2743 19431
rect 2685 19391 2743 19397
rect 2869 19431 2927 19437
rect 2869 19397 2881 19431
rect 2915 19428 2927 19431
rect 5718 19428 5724 19440
rect 2915 19400 5724 19428
rect 2915 19397 2927 19400
rect 2869 19391 2927 19397
rect 1486 19320 1492 19372
rect 1544 19360 1550 19372
rect 1762 19360 1768 19372
rect 1544 19332 1768 19360
rect 1544 19320 1550 19332
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 2038 19320 2044 19372
rect 2096 19320 2102 19372
rect 2130 19320 2136 19372
rect 2188 19320 2194 19372
rect 2222 19320 2228 19372
rect 2280 19360 2286 19372
rect 2884 19360 2912 19391
rect 5718 19388 5724 19400
rect 5776 19388 5782 19440
rect 2280 19332 2912 19360
rect 2961 19363 3019 19369
rect 2280 19320 2286 19332
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 4798 19360 4804 19372
rect 3007 19332 4804 19360
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 1581 19295 1639 19301
rect 1581 19261 1593 19295
rect 1627 19292 1639 19295
rect 1946 19292 1952 19304
rect 1627 19264 1952 19292
rect 1627 19261 1639 19264
rect 1581 19255 1639 19261
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 1104 19066 18860 19088
rect 1104 19014 3169 19066
rect 3221 19014 3233 19066
rect 3285 19014 3297 19066
rect 3349 19014 3361 19066
rect 3413 19014 3425 19066
rect 3477 19014 7608 19066
rect 7660 19014 7672 19066
rect 7724 19014 7736 19066
rect 7788 19014 7800 19066
rect 7852 19014 7864 19066
rect 7916 19014 12047 19066
rect 12099 19014 12111 19066
rect 12163 19014 12175 19066
rect 12227 19014 12239 19066
rect 12291 19014 12303 19066
rect 12355 19014 16486 19066
rect 16538 19014 16550 19066
rect 16602 19014 16614 19066
rect 16666 19014 16678 19066
rect 16730 19014 16742 19066
rect 16794 19014 18860 19066
rect 1104 18992 18860 19014
rect 3050 18912 3056 18964
rect 3108 18952 3114 18964
rect 3145 18955 3203 18961
rect 3145 18952 3157 18955
rect 3108 18924 3157 18952
rect 3108 18912 3114 18924
rect 3145 18921 3157 18924
rect 3191 18952 3203 18955
rect 3329 18955 3387 18961
rect 3191 18924 3280 18952
rect 3191 18921 3203 18924
rect 3145 18915 3203 18921
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 2961 18819 3019 18825
rect 2961 18816 2973 18819
rect 2832 18788 2973 18816
rect 2832 18776 2838 18788
rect 2961 18785 2973 18788
rect 3007 18785 3019 18819
rect 2961 18779 3019 18785
rect 3252 18760 3280 18924
rect 3329 18921 3341 18955
rect 3375 18952 3387 18955
rect 3786 18952 3792 18964
rect 3375 18924 3792 18952
rect 3375 18921 3387 18924
rect 3329 18915 3387 18921
rect 3786 18912 3792 18924
rect 3844 18912 3850 18964
rect 5905 18955 5963 18961
rect 5905 18921 5917 18955
rect 5951 18952 5963 18955
rect 6454 18952 6460 18964
rect 5951 18924 6460 18952
rect 5951 18921 5963 18924
rect 5905 18915 5963 18921
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 3145 18751 3203 18757
rect 3145 18748 3157 18751
rect 2372 18720 3157 18748
rect 2372 18708 2378 18720
rect 3145 18717 3157 18720
rect 3191 18717 3203 18751
rect 3145 18711 3203 18717
rect 3234 18708 3240 18760
rect 3292 18708 3298 18760
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18717 5043 18751
rect 4985 18711 5043 18717
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 5902 18748 5908 18760
rect 5399 18720 5908 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 2869 18683 2927 18689
rect 2869 18649 2881 18683
rect 2915 18680 2927 18683
rect 3602 18680 3608 18692
rect 2915 18652 3608 18680
rect 2915 18649 2927 18652
rect 2869 18643 2927 18649
rect 3602 18640 3608 18652
rect 3660 18640 3666 18692
rect 5000 18680 5028 18711
rect 5902 18708 5908 18720
rect 5960 18708 5966 18760
rect 6638 18680 6644 18692
rect 5000 18652 6644 18680
rect 6638 18640 6644 18652
rect 6696 18680 6702 18692
rect 6914 18680 6920 18692
rect 6696 18652 6920 18680
rect 6696 18640 6702 18652
rect 6914 18640 6920 18652
rect 6972 18640 6978 18692
rect 1104 18522 19019 18544
rect 1104 18470 5388 18522
rect 5440 18470 5452 18522
rect 5504 18470 5516 18522
rect 5568 18470 5580 18522
rect 5632 18470 5644 18522
rect 5696 18470 9827 18522
rect 9879 18470 9891 18522
rect 9943 18470 9955 18522
rect 10007 18470 10019 18522
rect 10071 18470 10083 18522
rect 10135 18470 14266 18522
rect 14318 18470 14330 18522
rect 14382 18470 14394 18522
rect 14446 18470 14458 18522
rect 14510 18470 14522 18522
rect 14574 18470 18705 18522
rect 18757 18470 18769 18522
rect 18821 18470 18833 18522
rect 18885 18470 18897 18522
rect 18949 18470 18961 18522
rect 19013 18470 19019 18522
rect 1104 18448 19019 18470
rect 2056 18312 3004 18340
rect 2056 18281 2084 18312
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 2976 18281 3004 18312
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2464 18244 2881 18272
rect 2464 18232 2470 18244
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18272 3019 18275
rect 3234 18272 3240 18284
rect 3007 18244 3240 18272
rect 3007 18241 3019 18244
rect 2961 18235 3019 18241
rect 3234 18232 3240 18244
rect 3292 18272 3298 18284
rect 4798 18272 4804 18284
rect 3292 18244 4804 18272
rect 3292 18232 3298 18244
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 2314 18204 2320 18216
rect 2271 18176 2320 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2314 18164 2320 18176
rect 2372 18204 2378 18216
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2372 18176 2789 18204
rect 2372 18164 2378 18176
rect 2777 18173 2789 18176
rect 2823 18173 2835 18207
rect 3053 18207 3111 18213
rect 3053 18204 3065 18207
rect 2777 18167 2835 18173
rect 2884 18176 3065 18204
rect 2884 18148 2912 18176
rect 3053 18173 3065 18176
rect 3099 18173 3111 18207
rect 3053 18167 3111 18173
rect 2866 18096 2872 18148
rect 2924 18096 2930 18148
rect 1857 18071 1915 18077
rect 1857 18037 1869 18071
rect 1903 18068 1915 18071
rect 2498 18068 2504 18080
rect 1903 18040 2504 18068
rect 1903 18037 1915 18040
rect 1857 18031 1915 18037
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 3050 18028 3056 18080
rect 3108 18068 3114 18080
rect 3237 18071 3295 18077
rect 3237 18068 3249 18071
rect 3108 18040 3249 18068
rect 3108 18028 3114 18040
rect 3237 18037 3249 18040
rect 3283 18037 3295 18071
rect 3237 18031 3295 18037
rect 1104 17978 18860 18000
rect 1104 17926 3169 17978
rect 3221 17926 3233 17978
rect 3285 17926 3297 17978
rect 3349 17926 3361 17978
rect 3413 17926 3425 17978
rect 3477 17926 7608 17978
rect 7660 17926 7672 17978
rect 7724 17926 7736 17978
rect 7788 17926 7800 17978
rect 7852 17926 7864 17978
rect 7916 17926 12047 17978
rect 12099 17926 12111 17978
rect 12163 17926 12175 17978
rect 12227 17926 12239 17978
rect 12291 17926 12303 17978
rect 12355 17926 16486 17978
rect 16538 17926 16550 17978
rect 16602 17926 16614 17978
rect 16666 17926 16678 17978
rect 16730 17926 16742 17978
rect 16794 17926 18860 17978
rect 1104 17904 18860 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 2590 17864 2596 17876
rect 1912 17836 2596 17864
rect 1912 17824 1918 17836
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 2958 17824 2964 17876
rect 3016 17824 3022 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 3510 17864 3516 17876
rect 3375 17836 3516 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17728 2191 17731
rect 3053 17731 3111 17737
rect 2179 17700 2728 17728
rect 2179 17697 2191 17700
rect 2133 17691 2191 17697
rect 2222 17620 2228 17672
rect 2280 17660 2286 17672
rect 2317 17663 2375 17669
rect 2317 17660 2329 17663
rect 2280 17632 2329 17660
rect 2280 17620 2286 17632
rect 2317 17629 2329 17632
rect 2363 17629 2375 17663
rect 2317 17623 2375 17629
rect 2406 17620 2412 17672
rect 2464 17620 2470 17672
rect 2130 17484 2136 17536
rect 2188 17484 2194 17536
rect 2590 17484 2596 17536
rect 2648 17524 2654 17536
rect 2700 17524 2728 17700
rect 3053 17697 3065 17731
rect 3099 17728 3111 17731
rect 3878 17728 3884 17740
rect 3099 17700 3884 17728
rect 3099 17697 3111 17700
rect 3053 17691 3111 17697
rect 3878 17688 3884 17700
rect 3936 17688 3942 17740
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 3510 17660 3516 17672
rect 3191 17632 3516 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 3510 17620 3516 17632
rect 3568 17620 3574 17672
rect 2869 17595 2927 17601
rect 2869 17561 2881 17595
rect 2915 17592 2927 17595
rect 3694 17592 3700 17604
rect 2915 17564 3700 17592
rect 2915 17561 2927 17564
rect 2869 17555 2927 17561
rect 3694 17552 3700 17564
rect 3752 17552 3758 17604
rect 3970 17524 3976 17536
rect 2648 17496 3976 17524
rect 2648 17484 2654 17496
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 1104 17434 19019 17456
rect 1104 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 5644 17434
rect 5696 17382 9827 17434
rect 9879 17382 9891 17434
rect 9943 17382 9955 17434
rect 10007 17382 10019 17434
rect 10071 17382 10083 17434
rect 10135 17382 14266 17434
rect 14318 17382 14330 17434
rect 14382 17382 14394 17434
rect 14446 17382 14458 17434
rect 14510 17382 14522 17434
rect 14574 17382 18705 17434
rect 18757 17382 18769 17434
rect 18821 17382 18833 17434
rect 18885 17382 18897 17434
rect 18949 17382 18961 17434
rect 19013 17382 19019 17434
rect 1104 17360 19019 17382
rect 2222 17144 2228 17196
rect 2280 17184 2286 17196
rect 2866 17184 2872 17196
rect 2280 17156 2872 17184
rect 2280 17144 2286 17156
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17184 3111 17187
rect 3786 17184 3792 17196
rect 3099 17156 3792 17184
rect 3099 17153 3111 17156
rect 3053 17147 3111 17153
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17184 3939 17187
rect 3970 17184 3976 17196
rect 3927 17156 3976 17184
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 2406 17116 2412 17128
rect 2004 17088 2412 17116
rect 2004 17076 2010 17088
rect 2406 17076 2412 17088
rect 2464 17116 2470 17128
rect 2685 17119 2743 17125
rect 2685 17116 2697 17119
rect 2464 17088 2697 17116
rect 2464 17076 2470 17088
rect 2685 17085 2697 17088
rect 2731 17085 2743 17119
rect 2685 17079 2743 17085
rect 4062 17076 4068 17128
rect 4120 17076 4126 17128
rect 2038 17008 2044 17060
rect 2096 17048 2102 17060
rect 3697 17051 3755 17057
rect 3697 17048 3709 17051
rect 2096 17020 3709 17048
rect 2096 17008 2102 17020
rect 3697 17017 3709 17020
rect 3743 17017 3755 17051
rect 3697 17011 3755 17017
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 7098 16980 7104 16992
rect 1728 16952 7104 16980
rect 1728 16940 1734 16952
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 1854 16736 1860 16788
rect 1912 16776 1918 16788
rect 7466 16776 7472 16788
rect 1912 16748 7472 16776
rect 1912 16736 1918 16748
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 2406 16668 2412 16720
rect 2464 16708 2470 16720
rect 2774 16708 2780 16720
rect 2464 16680 2780 16708
rect 2464 16668 2470 16680
rect 2774 16668 2780 16680
rect 2832 16668 2838 16720
rect 2958 16668 2964 16720
rect 3016 16668 3022 16720
rect 3234 16668 3240 16720
rect 3292 16708 3298 16720
rect 3786 16708 3792 16720
rect 3292 16680 3792 16708
rect 3292 16668 3298 16680
rect 3786 16668 3792 16680
rect 3844 16668 3850 16720
rect 934 16600 940 16652
rect 992 16640 998 16652
rect 1581 16643 1639 16649
rect 1581 16640 1593 16643
rect 992 16612 1593 16640
rect 992 16600 998 16612
rect 1581 16609 1593 16612
rect 1627 16609 1639 16643
rect 1581 16603 1639 16609
rect 2590 16600 2596 16652
rect 2648 16640 2654 16652
rect 3053 16643 3111 16649
rect 3053 16640 3065 16643
rect 2648 16612 3065 16640
rect 2648 16600 2654 16612
rect 3053 16609 3065 16612
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 3142 16600 3148 16652
rect 3200 16640 3206 16652
rect 3970 16640 3976 16652
rect 3200 16612 3976 16640
rect 3200 16600 3206 16612
rect 3970 16600 3976 16612
rect 4028 16600 4034 16652
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 5399 16612 5488 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 2869 16575 2927 16581
rect 2869 16541 2881 16575
rect 2915 16572 2927 16575
rect 3160 16572 3188 16600
rect 2915 16544 3188 16572
rect 5460 16572 5488 16612
rect 5810 16572 5816 16584
rect 5460 16544 5816 16572
rect 2915 16541 2927 16544
rect 2869 16535 2927 16541
rect 2792 16504 2820 16535
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 4062 16504 4068 16516
rect 2792 16476 4068 16504
rect 4062 16464 4068 16476
rect 4120 16464 4126 16516
rect 4982 16464 4988 16516
rect 5040 16504 5046 16516
rect 5086 16507 5144 16513
rect 5086 16504 5098 16507
rect 5040 16476 5098 16504
rect 5040 16464 5046 16476
rect 5086 16473 5098 16476
rect 5132 16473 5144 16507
rect 5086 16467 5144 16473
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3142 16436 3148 16448
rect 2832 16408 3148 16436
rect 2832 16396 2838 16408
rect 3142 16396 3148 16408
rect 3200 16396 3206 16448
rect 3602 16396 3608 16448
rect 3660 16436 3666 16448
rect 3973 16439 4031 16445
rect 3973 16436 3985 16439
rect 3660 16408 3985 16436
rect 3660 16396 3666 16408
rect 3973 16405 3985 16408
rect 4019 16405 4031 16439
rect 3973 16399 4031 16405
rect 1104 16346 19019 16368
rect 1104 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 5644 16346
rect 5696 16294 9827 16346
rect 9879 16294 9891 16346
rect 9943 16294 9955 16346
rect 10007 16294 10019 16346
rect 10071 16294 10083 16346
rect 10135 16294 14266 16346
rect 14318 16294 14330 16346
rect 14382 16294 14394 16346
rect 14446 16294 14458 16346
rect 14510 16294 14522 16346
rect 14574 16294 18705 16346
rect 18757 16294 18769 16346
rect 18821 16294 18833 16346
rect 18885 16294 18897 16346
rect 18949 16294 18961 16346
rect 19013 16294 19019 16346
rect 1104 16272 19019 16294
rect 1578 16192 1584 16244
rect 1636 16192 1642 16244
rect 1673 16235 1731 16241
rect 1673 16201 1685 16235
rect 1719 16232 1731 16235
rect 2406 16232 2412 16244
rect 1719 16204 2412 16232
rect 1719 16201 1731 16204
rect 1673 16195 1731 16201
rect 2406 16192 2412 16204
rect 2464 16192 2470 16244
rect 2682 16192 2688 16244
rect 2740 16232 2746 16244
rect 5169 16235 5227 16241
rect 2740 16204 4844 16232
rect 2740 16192 2746 16204
rect 1596 16164 1624 16192
rect 4034 16167 4092 16173
rect 4034 16164 4046 16167
rect 1596 16136 4046 16164
rect 4034 16133 4046 16136
rect 4080 16133 4092 16167
rect 4816 16164 4844 16204
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 5258 16232 5264 16244
rect 5215 16204 5264 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6178 16192 6184 16244
rect 6236 16232 6242 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 6236 16204 7941 16232
rect 6236 16192 6242 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 6794 16167 6852 16173
rect 6794 16164 6806 16167
rect 4816 16136 6806 16164
rect 4034 16127 4092 16133
rect 6794 16133 6806 16136
rect 6840 16133 6852 16167
rect 6794 16127 6852 16133
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 1762 16096 1768 16108
rect 1627 16068 1768 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 750 15920 756 15972
rect 808 15960 814 15972
rect 1872 15960 1900 16059
rect 2130 16056 2136 16108
rect 2188 16096 2194 16108
rect 2777 16099 2835 16105
rect 2777 16096 2789 16099
rect 2188 16068 2789 16096
rect 2188 16056 2194 16068
rect 2777 16065 2789 16068
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16096 3019 16099
rect 3142 16096 3148 16108
rect 3007 16068 3148 16096
rect 3007 16065 3019 16068
rect 2961 16059 3019 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 6270 16096 6276 16108
rect 3712 16068 6276 16096
rect 2590 15988 2596 16040
rect 2648 16028 2654 16040
rect 3712 16028 3740 16068
rect 6270 16056 6276 16068
rect 6328 16056 6334 16108
rect 2648 16000 3740 16028
rect 2648 15988 2654 16000
rect 3786 15988 3792 16040
rect 3844 15988 3850 16040
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 6549 16031 6607 16037
rect 6549 16028 6561 16031
rect 6236 16000 6561 16028
rect 6236 15988 6242 16000
rect 6549 15997 6561 16000
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 2682 15960 2688 15972
rect 808 15932 2688 15960
rect 808 15920 814 15932
rect 2682 15920 2688 15932
rect 2740 15960 2746 15972
rect 2866 15960 2872 15972
rect 2740 15932 2872 15960
rect 2740 15920 2746 15932
rect 2866 15920 2872 15932
rect 2924 15920 2930 15972
rect 6454 15960 6460 15972
rect 5092 15932 6460 15960
rect 1946 15852 1952 15904
rect 2004 15892 2010 15904
rect 2041 15895 2099 15901
rect 2041 15892 2053 15895
rect 2004 15864 2053 15892
rect 2004 15852 2010 15864
rect 2041 15861 2053 15864
rect 2087 15861 2099 15895
rect 2041 15855 2099 15861
rect 2130 15852 2136 15904
rect 2188 15892 2194 15904
rect 2590 15892 2596 15904
rect 2188 15864 2596 15892
rect 2188 15852 2194 15864
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 5092 15892 5120 15932
rect 6454 15920 6460 15932
rect 6512 15920 6518 15972
rect 2823 15864 5120 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 2130 15688 2136 15700
rect 1995 15660 2136 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2682 15648 2688 15700
rect 2740 15688 2746 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 2740 15660 2789 15688
rect 2740 15648 2746 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 2777 15651 2835 15657
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7524 15660 7849 15688
rect 7524 15648 7530 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15620 1639 15623
rect 2590 15620 2596 15632
rect 1627 15592 2596 15620
rect 1627 15589 1639 15592
rect 1581 15583 1639 15589
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 4617 15623 4675 15629
rect 4617 15620 4629 15623
rect 2746 15592 4629 15620
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 2746 15484 2774 15592
rect 4617 15589 4629 15592
rect 4663 15589 4675 15623
rect 4617 15583 4675 15589
rect 1452 15456 2774 15484
rect 1452 15444 1458 15456
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 4764 15456 5856 15484
rect 4764 15444 4770 15456
rect 1946 15376 1952 15428
rect 2004 15376 2010 15428
rect 2745 15419 2803 15425
rect 2745 15416 2757 15419
rect 2056 15388 2757 15416
rect 1762 15308 1768 15360
rect 1820 15348 1826 15360
rect 2056 15348 2084 15388
rect 2745 15385 2757 15388
rect 2791 15385 2803 15419
rect 2745 15379 2803 15385
rect 2866 15376 2872 15428
rect 2924 15416 2930 15428
rect 2961 15419 3019 15425
rect 2961 15416 2973 15419
rect 2924 15388 2973 15416
rect 2924 15376 2930 15388
rect 2961 15385 2973 15388
rect 3007 15385 3019 15419
rect 2961 15379 3019 15385
rect 5730 15419 5788 15425
rect 5730 15385 5742 15419
rect 5776 15385 5788 15419
rect 5828 15416 5856 15456
rect 5902 15444 5908 15496
rect 5960 15484 5966 15496
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 5960 15456 6009 15484
rect 5960 15444 5966 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 6457 15487 6515 15493
rect 6457 15484 6469 15487
rect 6236 15456 6469 15484
rect 6236 15444 6242 15456
rect 6457 15453 6469 15456
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 6702 15419 6760 15425
rect 6702 15416 6714 15419
rect 5828 15388 6714 15416
rect 5730 15379 5788 15385
rect 6702 15385 6714 15388
rect 6748 15385 6760 15419
rect 6702 15379 6760 15385
rect 1820 15320 2084 15348
rect 2133 15351 2191 15357
rect 1820 15308 1826 15320
rect 2133 15317 2145 15351
rect 2179 15348 2191 15351
rect 5074 15348 5080 15360
rect 2179 15320 5080 15348
rect 2179 15317 2191 15320
rect 2133 15311 2191 15317
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 5736 15348 5764 15379
rect 8846 15348 8852 15360
rect 5736 15320 8852 15348
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 1104 15258 19019 15280
rect 1104 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 5644 15258
rect 5696 15206 9827 15258
rect 9879 15206 9891 15258
rect 9943 15206 9955 15258
rect 10007 15206 10019 15258
rect 10071 15206 10083 15258
rect 10135 15206 14266 15258
rect 14318 15206 14330 15258
rect 14382 15206 14394 15258
rect 14446 15206 14458 15258
rect 14510 15206 14522 15258
rect 14574 15206 18705 15258
rect 18757 15206 18769 15258
rect 18821 15206 18833 15258
rect 18885 15206 18897 15258
rect 18949 15206 18961 15258
rect 19013 15206 19019 15258
rect 1104 15184 19019 15206
rect 2314 15104 2320 15156
rect 2372 15104 2378 15156
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 2866 15144 2872 15156
rect 2464 15116 2872 15144
rect 2464 15104 2470 15116
rect 2866 15104 2872 15116
rect 2924 15144 2930 15156
rect 4249 15147 4307 15153
rect 4249 15144 4261 15147
rect 2924 15116 4261 15144
rect 2924 15104 2930 15116
rect 4249 15113 4261 15116
rect 4295 15113 4307 15147
rect 4249 15107 4307 15113
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5902 15144 5908 15156
rect 5776 15116 5908 15144
rect 5776 15104 5782 15116
rect 5902 15104 5908 15116
rect 5960 15104 5966 15156
rect 7929 15147 7987 15153
rect 7929 15113 7941 15147
rect 7975 15144 7987 15147
rect 8110 15144 8116 15156
rect 7975 15116 8116 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 6822 15085 6828 15088
rect 6816 15076 6828 15085
rect 6783 15048 6828 15076
rect 6816 15039 6828 15048
rect 6822 15036 6828 15039
rect 6880 15036 6886 15088
rect 2682 14968 2688 15020
rect 2740 15008 2746 15020
rect 3430 15011 3488 15017
rect 3430 15008 3442 15011
rect 2740 14980 3442 15008
rect 2740 14968 2746 14980
rect 3430 14977 3442 14980
rect 3476 14977 3488 15011
rect 3430 14971 3488 14977
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 15008 5595 15011
rect 6270 15008 6276 15020
rect 5583 14980 6276 15008
rect 5583 14977 5595 14980
rect 5537 14971 5595 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 7926 14968 7932 15020
rect 7984 15008 7990 15020
rect 8110 15008 8116 15020
rect 7984 14980 8116 15008
rect 7984 14968 7990 14980
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 3697 14943 3755 14949
rect 3697 14909 3709 14943
rect 3743 14940 3755 14943
rect 3786 14940 3792 14952
rect 3743 14912 3792 14940
rect 3743 14909 3755 14912
rect 3697 14903 3755 14909
rect 3786 14900 3792 14912
rect 3844 14940 3850 14952
rect 3970 14940 3976 14952
rect 3844 14912 3976 14940
rect 3844 14900 3850 14912
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 5810 14900 5816 14952
rect 5868 14900 5874 14952
rect 6178 14900 6184 14952
rect 6236 14940 6242 14952
rect 6549 14943 6607 14949
rect 6549 14940 6561 14943
rect 6236 14912 6561 14940
rect 6236 14900 6242 14912
rect 6549 14909 6561 14912
rect 6595 14909 6607 14943
rect 6549 14903 6607 14909
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 4120 14572 4169 14600
rect 4120 14560 4126 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 4157 14563 4215 14569
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 5718 14600 5724 14612
rect 4304 14572 5724 14600
rect 4304 14560 4310 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 3418 14396 3424 14408
rect 2188 14368 3424 14396
rect 2188 14356 2194 14368
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 3970 14356 3976 14408
rect 4028 14396 4034 14408
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 4028 14368 5549 14396
rect 4028 14356 4034 14368
rect 5537 14365 5549 14368
rect 5583 14396 5595 14399
rect 5810 14396 5816 14408
rect 5583 14368 5816 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 6178 14356 6184 14408
rect 6236 14356 6242 14408
rect 6454 14405 6460 14408
rect 6448 14396 6460 14405
rect 6415 14368 6460 14396
rect 6448 14359 6460 14368
rect 6454 14356 6460 14359
rect 6512 14356 6518 14408
rect 1946 14288 1952 14340
rect 2004 14328 2010 14340
rect 2004 14300 5212 14328
rect 2004 14288 2010 14300
rect 5184 14260 5212 14300
rect 5258 14288 5264 14340
rect 5316 14337 5322 14340
rect 5316 14291 5328 14337
rect 5316 14288 5322 14291
rect 7561 14263 7619 14269
rect 7561 14260 7573 14263
rect 5184 14232 7573 14260
rect 7561 14229 7573 14232
rect 7607 14229 7619 14263
rect 7561 14223 7619 14229
rect 1104 14170 19019 14192
rect 1104 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 5644 14170
rect 5696 14118 9827 14170
rect 9879 14118 9891 14170
rect 9943 14118 9955 14170
rect 10007 14118 10019 14170
rect 10071 14118 10083 14170
rect 10135 14118 14266 14170
rect 14318 14118 14330 14170
rect 14382 14118 14394 14170
rect 14446 14118 14458 14170
rect 14510 14118 14522 14170
rect 14574 14118 18705 14170
rect 18757 14118 18769 14170
rect 18821 14118 18833 14170
rect 18885 14118 18897 14170
rect 18949 14118 18961 14170
rect 19013 14118 19019 14170
rect 1104 14096 19019 14118
rect 2682 14065 2688 14068
rect 2678 14056 2688 14065
rect 2643 14028 2688 14056
rect 2678 14019 2688 14028
rect 2682 14016 2688 14019
rect 2740 14016 2746 14068
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 5258 14056 5264 14068
rect 4764 14028 5264 14056
rect 4764 14016 4770 14028
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 5721 14059 5779 14065
rect 5721 14025 5733 14059
rect 5767 14056 5779 14059
rect 5902 14056 5908 14068
rect 5767 14028 5908 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 7929 14059 7987 14065
rect 7929 14025 7941 14059
rect 7975 14025 7987 14059
rect 7929 14019 7987 14025
rect 2777 13991 2835 13997
rect 2777 13957 2789 13991
rect 2823 13988 2835 13991
rect 3329 13991 3387 13997
rect 3329 13988 3341 13991
rect 2823 13960 3341 13988
rect 2823 13957 2835 13960
rect 2777 13951 2835 13957
rect 3329 13957 3341 13960
rect 3375 13957 3387 13991
rect 7944 13988 7972 14019
rect 3329 13951 3387 13957
rect 3896 13960 7972 13988
rect 1854 13880 1860 13932
rect 1912 13920 1918 13932
rect 2498 13920 2504 13932
rect 1912 13892 2504 13920
rect 1912 13880 1918 13892
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2866 13920 2872 13932
rect 2639 13892 2872 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 3050 13880 3056 13932
rect 3108 13920 3114 13932
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 3108 13892 3249 13920
rect 3108 13880 3114 13892
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 3418 13880 3424 13932
rect 3476 13880 3482 13932
rect 1210 13812 1216 13864
rect 1268 13852 1274 13864
rect 3896 13852 3924 13960
rect 4430 13880 4436 13932
rect 4488 13920 4494 13932
rect 4597 13923 4655 13929
rect 4597 13920 4609 13923
rect 4488 13892 4609 13920
rect 4488 13880 4494 13892
rect 4597 13889 4609 13892
rect 4643 13889 4655 13923
rect 4597 13883 4655 13889
rect 6816 13923 6874 13929
rect 6816 13889 6828 13923
rect 6862 13920 6874 13923
rect 8754 13920 8760 13932
rect 6862 13892 8760 13920
rect 6862 13889 6874 13892
rect 6816 13883 6874 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 1268 13824 3924 13852
rect 1268 13812 1274 13824
rect 3970 13812 3976 13864
rect 4028 13852 4034 13864
rect 4341 13855 4399 13861
rect 4341 13852 4353 13855
rect 4028 13824 4353 13852
rect 4028 13812 4034 13824
rect 4341 13821 4353 13824
rect 4387 13821 4399 13855
rect 4341 13815 4399 13821
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 6454 13852 6460 13864
rect 6236 13824 6460 13852
rect 6236 13812 6242 13824
rect 6454 13812 6460 13824
rect 6512 13852 6518 13864
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 6512 13824 6561 13852
rect 6512 13812 6518 13824
rect 6549 13821 6561 13824
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 2685 13515 2743 13521
rect 2685 13481 2697 13515
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 2961 13515 3019 13521
rect 2961 13481 2973 13515
rect 3007 13512 3019 13515
rect 4890 13512 4896 13524
rect 3007 13484 4896 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 2700 13444 2728 13475
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 3050 13444 3056 13456
rect 2700 13416 3056 13444
rect 3050 13404 3056 13416
rect 3108 13444 3114 13456
rect 4062 13444 4068 13456
rect 3108 13416 4068 13444
rect 3108 13404 3114 13416
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2406 13376 2412 13388
rect 2004 13348 2412 13376
rect 2004 13336 2010 13348
rect 2406 13336 2412 13348
rect 2464 13376 2470 13388
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 2464 13348 2605 13376
rect 2464 13336 2470 13348
rect 2593 13345 2605 13348
rect 2639 13345 2651 13379
rect 2593 13339 2651 13345
rect 2774 13268 2780 13320
rect 2832 13268 2838 13320
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 2866 13240 2872 13252
rect 2547 13212 2872 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 2866 13200 2872 13212
rect 2924 13200 2930 13252
rect 5258 13200 5264 13252
rect 5316 13200 5322 13252
rect 6454 13132 6460 13184
rect 6512 13172 6518 13184
rect 6549 13175 6607 13181
rect 6549 13172 6561 13175
rect 6512 13144 6561 13172
rect 6512 13132 6518 13144
rect 6549 13141 6561 13144
rect 6595 13141 6607 13175
rect 6549 13135 6607 13141
rect 1104 13082 19019 13104
rect 1104 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 5644 13082
rect 5696 13030 9827 13082
rect 9879 13030 9891 13082
rect 9943 13030 9955 13082
rect 10007 13030 10019 13082
rect 10071 13030 10083 13082
rect 10135 13030 14266 13082
rect 14318 13030 14330 13082
rect 14382 13030 14394 13082
rect 14446 13030 14458 13082
rect 14510 13030 14522 13082
rect 14574 13030 18705 13082
rect 18757 13030 18769 13082
rect 18821 13030 18833 13082
rect 18885 13030 18897 13082
rect 18949 13030 18961 13082
rect 19013 13030 19019 13082
rect 1104 13008 19019 13030
rect 2130 12928 2136 12980
rect 2188 12928 2194 12980
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7156 12940 7941 12968
rect 7156 12928 7162 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 2148 12900 2176 12928
rect 1872 12872 2176 12900
rect 6816 12903 6874 12909
rect 1872 12773 1900 12872
rect 6816 12869 6828 12903
rect 6862 12900 6874 12903
rect 8662 12900 8668 12912
rect 6862 12872 8668 12900
rect 6862 12869 6874 12872
rect 6816 12863 6874 12869
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 2774 12832 2780 12844
rect 2179 12804 2780 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 2774 12792 2780 12804
rect 2832 12832 2838 12844
rect 4062 12832 4068 12844
rect 2832 12804 4068 12832
rect 2832 12792 2838 12804
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12832 4399 12835
rect 5258 12832 5264 12844
rect 4387 12804 5264 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12733 1915 12767
rect 1857 12727 1915 12733
rect 6454 12724 6460 12776
rect 6512 12764 6518 12776
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 6512 12736 6561 12764
rect 6512 12724 6518 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 2038 12656 2044 12708
rect 2096 12696 2102 12708
rect 3602 12696 3608 12708
rect 2096 12668 3608 12696
rect 2096 12656 2102 12668
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 1118 12588 1124 12640
rect 1176 12628 1182 12640
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1176 12600 1961 12628
rect 1176 12588 1182 12600
rect 1949 12597 1961 12600
rect 1995 12597 2007 12631
rect 1949 12591 2007 12597
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3970 12628 3976 12640
rect 3099 12600 3976 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3694 12424 3700 12436
rect 2924 12396 3700 12424
rect 2924 12384 2930 12396
rect 3694 12384 3700 12396
rect 3752 12424 3758 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 3752 12396 7941 12424
rect 3752 12384 3758 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 934 12316 940 12368
rect 992 12356 998 12368
rect 1581 12359 1639 12365
rect 1581 12356 1593 12359
rect 992 12328 1593 12356
rect 992 12316 998 12328
rect 1581 12325 1593 12328
rect 1627 12325 1639 12359
rect 1581 12319 1639 12325
rect 4430 12288 4436 12300
rect 1780 12260 4436 12288
rect 1780 12229 1808 12260
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 5629 12291 5687 12297
rect 5629 12257 5641 12291
rect 5675 12288 5687 12291
rect 5994 12288 6000 12300
rect 5675 12260 6000 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 5994 12248 6000 12260
rect 6052 12288 6058 12300
rect 6454 12288 6460 12300
rect 6052 12260 6460 12288
rect 6052 12248 6058 12260
rect 6454 12248 6460 12260
rect 6512 12288 6518 12300
rect 6549 12291 6607 12297
rect 6549 12288 6561 12291
rect 6512 12260 6561 12288
rect 6512 12248 6518 12260
rect 6549 12257 6561 12260
rect 6595 12257 6607 12291
rect 6549 12251 6607 12257
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2314 12220 2320 12232
rect 2004 12192 2320 12220
rect 2004 12180 2010 12192
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 1670 12112 1676 12164
rect 1728 12152 1734 12164
rect 2130 12152 2136 12164
rect 1728 12124 2136 12152
rect 1728 12112 1734 12124
rect 2130 12112 2136 12124
rect 2188 12152 2194 12164
rect 2424 12152 2452 12183
rect 2188 12124 2452 12152
rect 2188 12112 2194 12124
rect 1026 12044 1032 12096
rect 1084 12084 1090 12096
rect 2608 12084 2636 12183
rect 2682 12180 2688 12232
rect 2740 12180 2746 12232
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 2866 12220 2872 12232
rect 2823 12192 2872 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3053 12155 3111 12161
rect 3053 12121 3065 12155
rect 3099 12152 3111 12155
rect 5362 12155 5420 12161
rect 5362 12152 5374 12155
rect 3099 12124 5374 12152
rect 3099 12121 3111 12124
rect 3053 12115 3111 12121
rect 5362 12121 5374 12124
rect 5408 12121 5420 12155
rect 5362 12115 5420 12121
rect 6816 12155 6874 12161
rect 6816 12121 6828 12155
rect 6862 12121 6874 12155
rect 6816 12115 6874 12121
rect 1084 12056 2636 12084
rect 1084 12044 1090 12056
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3510 12084 3516 12096
rect 2924 12056 3516 12084
rect 2924 12044 2930 12056
rect 3510 12044 3516 12056
rect 3568 12084 3574 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 3568 12056 4261 12084
rect 3568 12044 3574 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6840 12084 6868 12115
rect 6788 12056 6868 12084
rect 6788 12044 6794 12056
rect 1104 11994 19019 12016
rect 1104 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 5644 11994
rect 5696 11942 9827 11994
rect 9879 11942 9891 11994
rect 9943 11942 9955 11994
rect 10007 11942 10019 11994
rect 10071 11942 10083 11994
rect 10135 11942 14266 11994
rect 14318 11942 14330 11994
rect 14382 11942 14394 11994
rect 14446 11942 14458 11994
rect 14510 11942 14522 11994
rect 14574 11942 18705 11994
rect 18757 11942 18769 11994
rect 18821 11942 18833 11994
rect 18885 11942 18897 11994
rect 18949 11942 18961 11994
rect 19013 11942 19019 11994
rect 1104 11920 19019 11942
rect 2225 11883 2283 11889
rect 2225 11849 2237 11883
rect 2271 11880 2283 11883
rect 2314 11880 2320 11892
rect 2271 11852 2320 11880
rect 2271 11849 2283 11852
rect 2225 11843 2283 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 4706 11880 4712 11892
rect 3099 11852 4712 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 1762 11772 1768 11824
rect 1820 11772 1826 11824
rect 1854 11772 1860 11824
rect 1912 11812 1918 11824
rect 2130 11812 2136 11824
rect 1912 11784 2136 11812
rect 1912 11772 1918 11784
rect 2130 11772 2136 11784
rect 2188 11772 2194 11824
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 4028 11784 5396 11812
rect 4028 11772 4034 11784
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 2317 11747 2375 11753
rect 2317 11744 2329 11747
rect 1360 11716 2329 11744
rect 1360 11704 1366 11716
rect 2317 11713 2329 11716
rect 2363 11744 2375 11747
rect 2774 11744 2780 11756
rect 2363 11716 2780 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 2958 11704 2964 11756
rect 3016 11704 3022 11756
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 3510 11744 3516 11756
rect 3191 11716 3516 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 5368 11753 5396 11784
rect 5086 11747 5144 11753
rect 5086 11744 5098 11747
rect 4396 11716 5098 11744
rect 4396 11704 4402 11716
rect 5086 11713 5098 11716
rect 5132 11713 5144 11747
rect 5086 11707 5144 11713
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 6454 11744 6460 11756
rect 5776 11716 6460 11744
rect 5776 11704 5782 11716
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 2501 11679 2559 11685
rect 2501 11676 2513 11679
rect 2464 11648 2513 11676
rect 2464 11636 2470 11648
rect 2501 11645 2513 11648
rect 2547 11645 2559 11679
rect 2501 11639 2559 11645
rect 3602 11568 3608 11620
rect 3660 11608 3666 11620
rect 3973 11611 4031 11617
rect 3973 11608 3985 11611
rect 3660 11580 3985 11608
rect 3660 11568 3666 11580
rect 3973 11577 3985 11580
rect 4019 11577 4031 11611
rect 3973 11571 4031 11577
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1762 11336 1768 11348
rect 1452 11308 1768 11336
rect 1452 11296 1458 11308
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 4120 11308 7389 11336
rect 4120 11296 4126 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 7377 11299 7435 11305
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11200 1639 11203
rect 1670 11200 1676 11212
rect 1627 11172 1676 11200
rect 1627 11169 1639 11172
rect 1581 11163 1639 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 1946 11132 1952 11144
rect 1903 11104 1952 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 1578 11024 1584 11076
rect 1636 11024 1642 11076
rect 3602 11024 3608 11076
rect 3660 11064 3666 11076
rect 6242 11067 6300 11073
rect 6242 11064 6254 11067
rect 3660 11036 6254 11064
rect 3660 11024 3666 11036
rect 6242 11033 6254 11036
rect 6288 11033 6300 11067
rect 6242 11027 6300 11033
rect 1104 10906 19019 10928
rect 1104 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 5644 10906
rect 5696 10854 9827 10906
rect 9879 10854 9891 10906
rect 9943 10854 9955 10906
rect 10007 10854 10019 10906
rect 10071 10854 10083 10906
rect 10135 10854 14266 10906
rect 14318 10854 14330 10906
rect 14382 10854 14394 10906
rect 14446 10854 14458 10906
rect 14510 10854 14522 10906
rect 14574 10854 18705 10906
rect 18757 10854 18769 10906
rect 18821 10854 18833 10906
rect 18885 10854 18897 10906
rect 18949 10854 18961 10906
rect 19013 10854 19019 10906
rect 1104 10832 19019 10854
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 6420 10764 7941 10792
rect 6420 10752 6426 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 7929 10755 7987 10761
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6052 10628 6561 10656
rect 6052 10616 6058 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 9030 10656 9036 10668
rect 6871 10628 9036 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 4672 10220 5365 10248
rect 4672 10208 4678 10220
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 5353 10211 5411 10217
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 7101 10183 7159 10189
rect 7101 10180 7113 10183
rect 5316 10152 7113 10180
rect 5316 10140 5322 10152
rect 7101 10149 7113 10152
rect 7147 10149 7159 10183
rect 7101 10143 7159 10149
rect 3970 10072 3976 10124
rect 4028 10072 4034 10124
rect 934 10004 940 10056
rect 992 10044 998 10056
rect 4246 10053 4252 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 992 10016 1593 10044
rect 992 10004 998 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 4240 10007 4252 10053
rect 4246 10004 4252 10007
rect 4304 10004 4310 10056
rect 5810 9936 5816 9988
rect 5868 9936 5874 9988
rect 1104 9818 19019 9840
rect 1104 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 5644 9818
rect 5696 9766 9827 9818
rect 9879 9766 9891 9818
rect 9943 9766 9955 9818
rect 10007 9766 10019 9818
rect 10071 9766 10083 9818
rect 10135 9766 14266 9818
rect 14318 9766 14330 9818
rect 14382 9766 14394 9818
rect 14446 9766 14458 9818
rect 14510 9766 14522 9818
rect 14574 9766 18705 9818
rect 18757 9766 18769 9818
rect 18821 9766 18833 9818
rect 18885 9766 18897 9818
rect 18949 9766 18961 9818
rect 19013 9766 19019 9818
rect 1104 9744 19019 9766
rect 1762 9596 1768 9648
rect 1820 9636 1826 9648
rect 1857 9639 1915 9645
rect 1857 9636 1869 9639
rect 1820 9608 1869 9636
rect 1820 9596 1826 9608
rect 1857 9605 1869 9608
rect 1903 9605 1915 9639
rect 1857 9599 1915 9605
rect 1946 9596 1952 9648
rect 2004 9636 2010 9648
rect 2057 9639 2115 9645
rect 2057 9636 2069 9639
rect 2004 9608 2069 9636
rect 2004 9596 2010 9608
rect 2057 9605 2069 9608
rect 2103 9605 2115 9639
rect 2057 9599 2115 9605
rect 6549 9639 6607 9645
rect 6549 9605 6561 9639
rect 6595 9636 6607 9639
rect 6638 9636 6644 9648
rect 6595 9608 6644 9636
rect 6595 9605 6607 9608
rect 6549 9599 6607 9605
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8018 9500 8024 9512
rect 7975 9472 8024 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8202 9460 8208 9512
rect 8260 9460 8266 9512
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2130 9364 2136 9376
rect 2087 9336 2136 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 4154 9364 4160 9376
rect 2271 9336 4160 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 3142 9120 3148 9172
rect 3200 9160 3206 9172
rect 3970 9160 3976 9172
rect 3200 9132 3976 9160
rect 3200 9120 3206 9132
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 1486 9052 1492 9104
rect 1544 9092 1550 9104
rect 1544 9064 4016 9092
rect 1544 9052 1550 9064
rect 3988 9036 4016 9064
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 9024 2007 9027
rect 2038 9024 2044 9036
rect 1995 8996 2044 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2038 8984 2044 8996
rect 2096 9024 2102 9036
rect 2498 9024 2504 9036
rect 2096 8996 2504 9024
rect 2096 8984 2102 8996
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 3970 8984 3976 9036
rect 4028 8984 4034 9036
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 1854 8956 1860 8968
rect 1627 8928 1860 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 1394 8848 1400 8900
rect 1452 8888 1458 8900
rect 1673 8891 1731 8897
rect 1673 8888 1685 8891
rect 1452 8860 1685 8888
rect 1452 8848 1458 8860
rect 1673 8857 1685 8860
rect 1719 8857 1731 8891
rect 1673 8851 1731 8857
rect 1780 8860 2636 8888
rect 1780 8829 1808 8860
rect 2608 8832 2636 8860
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8789 1823 8823
rect 1765 8783 1823 8789
rect 1946 8780 1952 8832
rect 2004 8780 2010 8832
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 3786 8820 3792 8832
rect 2648 8792 3792 8820
rect 2648 8780 2654 8792
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 1104 8730 19019 8752
rect 1104 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 5644 8730
rect 5696 8678 9827 8730
rect 9879 8678 9891 8730
rect 9943 8678 9955 8730
rect 10007 8678 10019 8730
rect 10071 8678 10083 8730
rect 10135 8678 14266 8730
rect 14318 8678 14330 8730
rect 14382 8678 14394 8730
rect 14446 8678 14458 8730
rect 14510 8678 14522 8730
rect 14574 8678 18705 8730
rect 18757 8678 18769 8730
rect 18821 8678 18833 8730
rect 18885 8678 18897 8730
rect 18949 8678 18961 8730
rect 19013 8678 19019 8730
rect 1104 8656 19019 8678
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 2869 8619 2927 8625
rect 2869 8616 2881 8619
rect 2832 8588 2881 8616
rect 2832 8576 2838 8588
rect 2869 8585 2881 8588
rect 2915 8616 2927 8619
rect 3050 8616 3056 8628
rect 2915 8588 3056 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 4856 8588 5181 8616
rect 4856 8576 4862 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 2682 8508 2688 8560
rect 2740 8508 2746 8560
rect 4056 8551 4114 8557
rect 4056 8517 4068 8551
rect 4102 8548 4114 8551
rect 6546 8548 6552 8560
rect 4102 8520 6552 8548
rect 4102 8517 4114 8520
rect 4056 8511 4114 8517
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8480 2835 8483
rect 2958 8480 2964 8492
rect 2823 8452 2964 8480
rect 2823 8449 2835 8452
rect 2777 8443 2835 8449
rect 2958 8440 2964 8452
rect 3016 8480 3022 8492
rect 3694 8480 3700 8492
rect 3016 8452 3700 8480
rect 3016 8440 3022 8452
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 2314 8372 2320 8424
rect 2372 8372 2378 8424
rect 3050 8372 3056 8424
rect 3108 8372 3114 8424
rect 3786 8372 3792 8424
rect 3844 8372 3850 8424
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 2866 7936 2872 7948
rect 2363 7908 2872 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 750 7828 756 7880
rect 808 7868 814 7880
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 808 7840 2145 7868
rect 808 7828 814 7840
rect 2133 7837 2145 7840
rect 2179 7868 2191 7871
rect 3694 7868 3700 7880
rect 2179 7840 3700 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 1949 7735 2007 7741
rect 1949 7732 1961 7735
rect 1912 7704 1961 7732
rect 1912 7692 1918 7704
rect 1949 7701 1961 7704
rect 1995 7701 2007 7735
rect 1949 7695 2007 7701
rect 1104 7642 19019 7664
rect 1104 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 5644 7642
rect 5696 7590 9827 7642
rect 9879 7590 9891 7642
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7590 10083 7642
rect 10135 7590 14266 7642
rect 14318 7590 14330 7642
rect 14382 7590 14394 7642
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7590 18705 7642
rect 18757 7590 18769 7642
rect 18821 7590 18833 7642
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 7190 7528 7196 7540
rect 6687 7500 7196 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 1302 7420 1308 7472
rect 1360 7460 1366 7472
rect 7776 7463 7834 7469
rect 1360 7432 2544 7460
rect 1360 7420 1366 7432
rect 2222 7352 2228 7404
rect 2280 7352 2286 7404
rect 2406 7352 2412 7404
rect 2464 7352 2470 7404
rect 2516 7401 2544 7432
rect 7776 7429 7788 7463
rect 7822 7460 7834 7463
rect 8386 7460 8392 7472
rect 7822 7432 8392 7460
rect 7822 7429 7834 7432
rect 7776 7423 7834 7429
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8202 7392 8208 7404
rect 8067 7364 8208 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 2314 7284 2320 7336
rect 2372 7284 2378 7336
rect 2038 7148 2044 7200
rect 2096 7148 2102 7200
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 6270 6984 6276 6996
rect 1719 6956 6276 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 1854 6876 1860 6928
rect 1912 6916 1918 6928
rect 1912 6888 2268 6916
rect 1912 6876 1918 6888
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 1452 6820 1992 6848
rect 1452 6808 1458 6820
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1964 6789 1992 6820
rect 2240 6792 2268 6888
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 2556 6820 2789 6848
rect 2556 6808 2562 6820
rect 2777 6817 2789 6820
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3844 6820 3985 6848
rect 3844 6808 3850 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1636 6752 1685 6780
rect 1636 6740 1642 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 1995 6752 2176 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 1857 6715 1915 6721
rect 1857 6712 1869 6715
rect 1688 6684 1869 6712
rect 1688 6656 1716 6684
rect 1857 6681 1869 6684
rect 1903 6681 1915 6715
rect 1857 6675 1915 6681
rect 1670 6604 1676 6656
rect 1728 6604 1734 6656
rect 2148 6644 2176 6752
rect 2222 6740 2228 6792
rect 2280 6780 2286 6792
rect 2409 6783 2467 6789
rect 2409 6780 2421 6783
rect 2280 6752 2421 6780
rect 2280 6740 2286 6752
rect 2409 6749 2421 6752
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 2958 6780 2964 6792
rect 2915 6752 2964 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 2958 6740 2964 6752
rect 3016 6780 3022 6792
rect 3878 6780 3884 6792
rect 3016 6752 3884 6780
rect 3016 6740 3022 6752
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4240 6783 4298 6789
rect 4240 6749 4252 6783
rect 4286 6780 4298 6783
rect 5166 6780 5172 6792
rect 4286 6752 5172 6780
rect 4286 6749 4298 6752
rect 4240 6743 4298 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 7098 6672 7104 6724
rect 7156 6712 7162 6724
rect 8202 6712 8208 6724
rect 7156 6684 8208 6712
rect 7156 6672 7162 6684
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 2148 6616 2513 6644
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 2682 6604 2688 6656
rect 2740 6604 2746 6656
rect 3050 6604 3056 6656
rect 3108 6604 3114 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 5353 6647 5411 6653
rect 5353 6644 5365 6647
rect 4028 6616 5365 6644
rect 4028 6604 4034 6616
rect 5353 6613 5365 6616
rect 5399 6613 5411 6647
rect 5353 6607 5411 6613
rect 1104 6554 19019 6576
rect 1104 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 5644 6554
rect 5696 6502 9827 6554
rect 9879 6502 9891 6554
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6502 10083 6554
rect 10135 6502 14266 6554
rect 14318 6502 14330 6554
rect 14382 6502 14394 6554
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6502 18705 6554
rect 18757 6502 18769 6554
rect 18821 6502 18833 6554
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 2498 6440 2504 6452
rect 1728 6412 2504 6440
rect 1728 6400 1734 6412
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 4614 6400 4620 6452
rect 4672 6400 4678 6452
rect 6288 6412 7236 6440
rect 3050 6372 3056 6384
rect 2240 6344 3056 6372
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 2240 6313 2268 6344
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 5752 6375 5810 6381
rect 5752 6341 5764 6375
rect 5798 6372 5810 6375
rect 6288 6372 6316 6412
rect 7098 6372 7104 6384
rect 5798 6344 6316 6372
rect 6564 6344 7104 6372
rect 5798 6341 5810 6344
rect 5752 6335 5810 6341
rect 6564 6316 6592 6344
rect 7098 6332 7104 6344
rect 7156 6332 7162 6384
rect 2041 6307 2099 6313
rect 2041 6304 2053 6307
rect 1912 6276 2053 6304
rect 1912 6264 1918 6276
rect 2041 6273 2053 6276
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 2332 6236 2360 6267
rect 2406 6264 2412 6316
rect 2464 6264 2470 6316
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 6546 6304 6552 6316
rect 6043 6276 6552 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6822 6313 6828 6316
rect 6816 6267 6828 6313
rect 6822 6264 6828 6267
rect 6880 6264 6886 6316
rect 7208 6304 7236 6412
rect 7282 6400 7288 6452
rect 7340 6440 7346 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7340 6412 7941 6440
rect 7340 6400 7346 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 9674 6304 9680 6316
rect 7208 6276 9680 6304
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 2004 6208 2360 6236
rect 2004 6196 2010 6208
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6100 2743 6103
rect 4890 6100 4896 6112
rect 2731 6072 4896 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 2501 5899 2559 5905
rect 2501 5896 2513 5899
rect 2464 5868 2513 5896
rect 2464 5856 2470 5868
rect 2501 5865 2513 5868
rect 2547 5865 2559 5899
rect 2501 5859 2559 5865
rect 6546 5856 6552 5908
rect 6604 5856 6610 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 8478 5896 8484 5908
rect 6880 5868 8484 5896
rect 6880 5856 6886 5868
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2958 5692 2964 5704
rect 2639 5664 2964 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 934 5584 940 5636
rect 992 5624 998 5636
rect 1581 5627 1639 5633
rect 1581 5624 1593 5627
rect 992 5596 1593 5624
rect 992 5584 998 5596
rect 1581 5593 1593 5596
rect 1627 5593 1639 5627
rect 1581 5587 1639 5593
rect 1762 5584 1768 5636
rect 1820 5584 1826 5636
rect 1104 5466 19019 5488
rect 1104 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 5644 5466
rect 5696 5414 9827 5466
rect 9879 5414 9891 5466
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5414 10083 5466
rect 10135 5414 14266 5466
rect 14318 5414 14330 5466
rect 14382 5414 14394 5466
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5414 18705 5466
rect 18757 5414 18769 5466
rect 18821 5414 18833 5466
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 2038 5352 2044 5364
rect 1995 5324 2044 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3786 5352 3792 5364
rect 3099 5324 3792 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8110 5352 8116 5364
rect 7975 5324 8116 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 5258 5284 5264 5296
rect 4387 5256 5264 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 6816 5287 6874 5293
rect 6816 5253 6828 5287
rect 6862 5284 6874 5287
rect 8570 5284 8576 5296
rect 6862 5256 8576 5284
rect 6862 5253 6874 5256
rect 6816 5247 6874 5253
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 1394 5176 1400 5228
rect 1452 5216 1458 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1452 5188 1593 5216
rect 1452 5176 1458 5188
rect 1581 5185 1593 5188
rect 1627 5216 1639 5219
rect 1854 5216 1860 5228
rect 1627 5188 1860 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2038 5176 2044 5228
rect 2096 5216 2102 5228
rect 3602 5216 3608 5228
rect 2096 5188 3608 5216
rect 2096 5176 2102 5188
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 2133 5083 2191 5089
rect 2133 5049 2145 5083
rect 2179 5080 2191 5083
rect 4982 5080 4988 5092
rect 2179 5052 4988 5080
rect 2179 5049 2191 5052
rect 2133 5043 2191 5049
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 1946 4972 1952 5024
rect 2004 4972 2010 5024
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 2041 4811 2099 4817
rect 2041 4808 2053 4811
rect 1820 4780 2053 4808
rect 1820 4768 1826 4780
rect 2041 4777 2053 4780
rect 2087 4777 2099 4811
rect 6546 4808 6552 4820
rect 2041 4771 2099 4777
rect 6196 4780 6552 4808
rect 3421 4675 3479 4681
rect 3421 4641 3433 4675
rect 3467 4672 3479 4675
rect 3786 4672 3792 4684
rect 3467 4644 3792 4672
rect 3467 4641 3479 4644
rect 3421 4635 3479 4641
rect 3786 4632 3792 4644
rect 3844 4672 3850 4684
rect 6196 4681 6224 4780
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 4249 4675 4307 4681
rect 4249 4672 4261 4675
rect 3844 4644 4261 4672
rect 3844 4632 3850 4644
rect 4249 4641 4261 4644
rect 4295 4641 4307 4675
rect 4249 4635 4307 4641
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 3165 4607 3223 4613
rect 3165 4573 3177 4607
rect 3211 4604 3223 4607
rect 4062 4604 4068 4616
rect 3211 4576 4068 4604
rect 3211 4573 3223 4576
rect 3165 4567 3223 4573
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4516 4607 4574 4613
rect 4516 4573 4528 4607
rect 4562 4604 4574 4607
rect 4798 4604 4804 4616
rect 4562 4576 4804 4604
rect 4562 4573 4574 4576
rect 4516 4567 4574 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 6454 4613 6460 4616
rect 6448 4567 6460 4613
rect 6454 4564 6460 4567
rect 6512 4564 6518 4616
rect 7374 4536 7380 4548
rect 5644 4508 7380 4536
rect 5644 4477 5672 4508
rect 7374 4496 7380 4508
rect 7432 4496 7438 4548
rect 5629 4471 5687 4477
rect 5629 4437 5641 4471
rect 5675 4437 5687 4471
rect 5629 4431 5687 4437
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 7561 4471 7619 4477
rect 7561 4468 7573 4471
rect 6052 4440 7573 4468
rect 6052 4428 6058 4440
rect 7561 4437 7573 4440
rect 7607 4437 7619 4471
rect 7561 4431 7619 4437
rect 1104 4378 19019 4400
rect 1104 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 5644 4378
rect 5696 4326 9827 4378
rect 9879 4326 9891 4378
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4326 10083 4378
rect 10135 4326 14266 4378
rect 14318 4326 14330 4378
rect 14382 4326 14394 4378
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4326 18705 4378
rect 18757 4326 18769 4378
rect 18821 4326 18833 4378
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 2700 4236 3004 4264
rect 1118 4156 1124 4208
rect 1176 4196 1182 4208
rect 1949 4199 2007 4205
rect 1949 4196 1961 4199
rect 1176 4168 1961 4196
rect 1176 4156 1182 4168
rect 1949 4165 1961 4168
rect 1995 4165 2007 4199
rect 2700 4196 2728 4236
rect 1949 4159 2007 4165
rect 2608 4168 2728 4196
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 2608 4128 2636 4168
rect 2774 4156 2780 4208
rect 2832 4156 2838 4208
rect 1765 4091 1823 4097
rect 2056 4100 2636 4128
rect 2685 4131 2743 4137
rect 1780 4060 1808 4091
rect 2056 4060 2084 4100
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2792 4128 2820 4156
rect 2731 4100 2820 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2866 4088 2872 4140
rect 2924 4088 2930 4140
rect 1780 4032 2084 4060
rect 2590 4020 2596 4072
rect 2648 4020 2654 4072
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2976 4060 3004 4236
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5178 4131 5236 4137
rect 5178 4128 5190 4131
rect 4948 4100 5190 4128
rect 4948 4088 4954 4100
rect 5178 4097 5190 4100
rect 5224 4097 5236 4131
rect 5178 4091 5236 4097
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 6270 4128 6276 4140
rect 5491 4100 6276 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 6270 4088 6276 4100
rect 6328 4128 6334 4140
rect 6546 4128 6552 4140
rect 6328 4100 6552 4128
rect 6328 4088 6334 4100
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 3050 4060 3056 4072
rect 2823 4032 3056 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 6086 4020 6092 4072
rect 6144 4060 6150 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 6144 4032 7941 4060
rect 6144 4020 6150 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 2038 3992 2044 4004
rect 1995 3964 2044 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 2038 3952 2044 3964
rect 2096 3952 2102 4004
rect 2958 3952 2964 4004
rect 3016 3992 3022 4004
rect 4065 3995 4123 4001
rect 4065 3992 4077 3995
rect 3016 3964 4077 3992
rect 3016 3952 3022 3964
rect 4065 3961 4077 3964
rect 4111 3961 4123 3995
rect 4065 3955 4123 3961
rect 2409 3927 2467 3933
rect 2409 3893 2421 3927
rect 2455 3924 2467 3927
rect 2590 3924 2596 3936
rect 2455 3896 2596 3924
rect 2455 3893 2467 3896
rect 2409 3887 2467 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2593 3723 2651 3729
rect 2593 3720 2605 3723
rect 2004 3692 2605 3720
rect 2004 3680 2010 3692
rect 2593 3689 2605 3692
rect 2639 3689 2651 3723
rect 2593 3683 2651 3689
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 6730 3720 6736 3732
rect 2823 3692 6736 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7837 3723 7895 3729
rect 7837 3689 7849 3723
rect 7883 3720 7895 3723
rect 9122 3720 9128 3732
rect 7883 3692 9128 3720
rect 7883 3689 7895 3692
rect 7837 3683 7895 3689
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 2225 3655 2283 3661
rect 2225 3621 2237 3655
rect 2271 3652 2283 3655
rect 2314 3652 2320 3664
rect 2271 3624 2320 3652
rect 2271 3621 2283 3624
rect 2225 3615 2283 3621
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 3510 3584 3516 3596
rect 1728 3556 3516 3584
rect 1728 3544 1734 3556
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 3786 3544 3792 3596
rect 3844 3584 3850 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 3844 3556 3985 3584
rect 3844 3544 3850 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 3973 3547 4031 3553
rect 6270 3544 6276 3596
rect 6328 3544 6334 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 7006 3584 7012 3596
rect 6595 3556 7012 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 4246 3525 4252 3528
rect 4240 3479 4252 3525
rect 4246 3476 4252 3479
rect 4304 3476 4310 3528
rect 4982 3476 4988 3528
rect 5040 3516 5046 3528
rect 5810 3516 5816 3528
rect 5040 3488 5816 3516
rect 5040 3476 5046 3488
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 2590 3408 2596 3460
rect 2648 3408 2654 3460
rect 842 3340 848 3392
rect 900 3380 906 3392
rect 5353 3383 5411 3389
rect 5353 3380 5365 3383
rect 900 3352 5365 3380
rect 900 3340 906 3352
rect 5353 3349 5365 3352
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 1104 3290 19019 3312
rect 1104 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 5644 3290
rect 5696 3238 9827 3290
rect 9879 3238 9891 3290
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3238 10083 3290
rect 10135 3238 14266 3290
rect 14318 3238 14330 3290
rect 14382 3238 14394 3290
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3238 18705 3290
rect 18757 3238 18769 3290
rect 18821 3238 18833 3290
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 2130 3136 2136 3188
rect 2188 3136 2194 3188
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4212 3148 4292 3176
rect 4212 3136 4218 3148
rect 4264 3117 4292 3148
rect 4240 3111 4298 3117
rect 4240 3077 4252 3111
rect 4286 3077 4298 3111
rect 4240 3071 4298 3077
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1636 3012 1961 3040
rect 1636 3000 1642 3012
rect 1949 3009 1961 3012
rect 1995 3040 2007 3043
rect 2222 3040 2228 3052
rect 1995 3012 2228 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3844 3012 3985 3040
rect 3844 3000 3850 3012
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 1688 2836 1716 2935
rect 1762 2932 1768 2984
rect 1820 2932 1826 2984
rect 1854 2932 1860 2984
rect 1912 2932 1918 2984
rect 2682 2836 2688 2848
rect 1688 2808 2688 2836
rect 2682 2796 2688 2808
rect 2740 2836 2746 2848
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 2740 2808 5365 2836
rect 2740 2796 2746 2808
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 5353 2799 5411 2805
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 1210 2592 1216 2644
rect 1268 2632 1274 2644
rect 1673 2635 1731 2641
rect 1673 2632 1685 2635
rect 1268 2604 1685 2632
rect 1268 2592 1274 2604
rect 1673 2601 1685 2604
rect 1719 2601 1731 2635
rect 1673 2595 1731 2601
rect 3694 2592 3700 2644
rect 3752 2632 3758 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 3752 2604 5365 2632
rect 3752 2592 3758 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 934 2456 940 2508
rect 992 2496 998 2508
rect 2317 2499 2375 2505
rect 2317 2496 2329 2499
rect 992 2468 2329 2496
rect 992 2456 998 2468
rect 2317 2465 2329 2468
rect 2363 2465 2375 2499
rect 2317 2459 2375 2465
rect 3786 2456 3792 2508
rect 3844 2496 3850 2508
rect 3973 2499 4031 2505
rect 3973 2496 3985 2499
rect 3844 2468 3985 2496
rect 3844 2456 3850 2468
rect 3973 2465 3985 2468
rect 4019 2465 4031 2499
rect 3973 2459 4031 2465
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 15381 2499 15439 2505
rect 15381 2496 15393 2499
rect 8996 2468 15393 2496
rect 8996 2456 9002 2468
rect 15381 2465 15393 2468
rect 15427 2465 15439 2499
rect 15381 2459 15439 2465
rect 1578 2388 1584 2440
rect 1636 2388 1642 2440
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 1780 2360 1808 2391
rect 1854 2388 1860 2440
rect 1912 2388 1918 2440
rect 4240 2431 4298 2437
rect 4240 2397 4252 2431
rect 4286 2428 4298 2431
rect 5074 2428 5080 2440
rect 4286 2400 5080 2428
rect 4286 2397 4298 2400
rect 4240 2391 4298 2397
rect 5074 2388 5080 2400
rect 5132 2388 5138 2440
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 1946 2360 1952 2372
rect 1780 2332 1952 2360
rect 1946 2320 1952 2332
rect 2004 2320 2010 2372
rect 1104 2202 19019 2224
rect 1104 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 5644 2202
rect 5696 2150 9827 2202
rect 9879 2150 9891 2202
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2150 10083 2202
rect 10135 2150 14266 2202
rect 14318 2150 14330 2202
rect 14382 2150 14394 2202
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2150 18705 2202
rect 18757 2150 18769 2202
rect 18821 2150 18833 2202
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
<< via1 >>
rect 3169 47302 3221 47354
rect 3233 47302 3285 47354
rect 3297 47302 3349 47354
rect 3361 47302 3413 47354
rect 3425 47302 3477 47354
rect 7608 47302 7660 47354
rect 7672 47302 7724 47354
rect 7736 47302 7788 47354
rect 7800 47302 7852 47354
rect 7864 47302 7916 47354
rect 12047 47302 12099 47354
rect 12111 47302 12163 47354
rect 12175 47302 12227 47354
rect 12239 47302 12291 47354
rect 12303 47302 12355 47354
rect 16486 47302 16538 47354
rect 16550 47302 16602 47354
rect 16614 47302 16666 47354
rect 16678 47302 16730 47354
rect 16742 47302 16794 47354
rect 940 47132 992 47184
rect 1400 46928 1452 46980
rect 5388 46758 5440 46810
rect 5452 46758 5504 46810
rect 5516 46758 5568 46810
rect 5580 46758 5632 46810
rect 5644 46758 5696 46810
rect 9827 46758 9879 46810
rect 9891 46758 9943 46810
rect 9955 46758 10007 46810
rect 10019 46758 10071 46810
rect 10083 46758 10135 46810
rect 14266 46758 14318 46810
rect 14330 46758 14382 46810
rect 14394 46758 14446 46810
rect 14458 46758 14510 46810
rect 14522 46758 14574 46810
rect 18705 46758 18757 46810
rect 18769 46758 18821 46810
rect 18833 46758 18885 46810
rect 18897 46758 18949 46810
rect 18961 46758 19013 46810
rect 3169 46214 3221 46266
rect 3233 46214 3285 46266
rect 3297 46214 3349 46266
rect 3361 46214 3413 46266
rect 3425 46214 3477 46266
rect 7608 46214 7660 46266
rect 7672 46214 7724 46266
rect 7736 46214 7788 46266
rect 7800 46214 7852 46266
rect 7864 46214 7916 46266
rect 12047 46214 12099 46266
rect 12111 46214 12163 46266
rect 12175 46214 12227 46266
rect 12239 46214 12291 46266
rect 12303 46214 12355 46266
rect 16486 46214 16538 46266
rect 16550 46214 16602 46266
rect 16614 46214 16666 46266
rect 16678 46214 16730 46266
rect 16742 46214 16794 46266
rect 5388 45670 5440 45722
rect 5452 45670 5504 45722
rect 5516 45670 5568 45722
rect 5580 45670 5632 45722
rect 5644 45670 5696 45722
rect 9827 45670 9879 45722
rect 9891 45670 9943 45722
rect 9955 45670 10007 45722
rect 10019 45670 10071 45722
rect 10083 45670 10135 45722
rect 14266 45670 14318 45722
rect 14330 45670 14382 45722
rect 14394 45670 14446 45722
rect 14458 45670 14510 45722
rect 14522 45670 14574 45722
rect 18705 45670 18757 45722
rect 18769 45670 18821 45722
rect 18833 45670 18885 45722
rect 18897 45670 18949 45722
rect 18961 45670 19013 45722
rect 3169 45126 3221 45178
rect 3233 45126 3285 45178
rect 3297 45126 3349 45178
rect 3361 45126 3413 45178
rect 3425 45126 3477 45178
rect 7608 45126 7660 45178
rect 7672 45126 7724 45178
rect 7736 45126 7788 45178
rect 7800 45126 7852 45178
rect 7864 45126 7916 45178
rect 12047 45126 12099 45178
rect 12111 45126 12163 45178
rect 12175 45126 12227 45178
rect 12239 45126 12291 45178
rect 12303 45126 12355 45178
rect 16486 45126 16538 45178
rect 16550 45126 16602 45178
rect 16614 45126 16666 45178
rect 16678 45126 16730 45178
rect 16742 45126 16794 45178
rect 940 44820 992 44872
rect 5388 44582 5440 44634
rect 5452 44582 5504 44634
rect 5516 44582 5568 44634
rect 5580 44582 5632 44634
rect 5644 44582 5696 44634
rect 9827 44582 9879 44634
rect 9891 44582 9943 44634
rect 9955 44582 10007 44634
rect 10019 44582 10071 44634
rect 10083 44582 10135 44634
rect 14266 44582 14318 44634
rect 14330 44582 14382 44634
rect 14394 44582 14446 44634
rect 14458 44582 14510 44634
rect 14522 44582 14574 44634
rect 18705 44582 18757 44634
rect 18769 44582 18821 44634
rect 18833 44582 18885 44634
rect 18897 44582 18949 44634
rect 18961 44582 19013 44634
rect 3169 44038 3221 44090
rect 3233 44038 3285 44090
rect 3297 44038 3349 44090
rect 3361 44038 3413 44090
rect 3425 44038 3477 44090
rect 7608 44038 7660 44090
rect 7672 44038 7724 44090
rect 7736 44038 7788 44090
rect 7800 44038 7852 44090
rect 7864 44038 7916 44090
rect 12047 44038 12099 44090
rect 12111 44038 12163 44090
rect 12175 44038 12227 44090
rect 12239 44038 12291 44090
rect 12303 44038 12355 44090
rect 16486 44038 16538 44090
rect 16550 44038 16602 44090
rect 16614 44038 16666 44090
rect 16678 44038 16730 44090
rect 16742 44038 16794 44090
rect 5388 43494 5440 43546
rect 5452 43494 5504 43546
rect 5516 43494 5568 43546
rect 5580 43494 5632 43546
rect 5644 43494 5696 43546
rect 9827 43494 9879 43546
rect 9891 43494 9943 43546
rect 9955 43494 10007 43546
rect 10019 43494 10071 43546
rect 10083 43494 10135 43546
rect 14266 43494 14318 43546
rect 14330 43494 14382 43546
rect 14394 43494 14446 43546
rect 14458 43494 14510 43546
rect 14522 43494 14574 43546
rect 18705 43494 18757 43546
rect 18769 43494 18821 43546
rect 18833 43494 18885 43546
rect 18897 43494 18949 43546
rect 18961 43494 19013 43546
rect 3169 42950 3221 43002
rect 3233 42950 3285 43002
rect 3297 42950 3349 43002
rect 3361 42950 3413 43002
rect 3425 42950 3477 43002
rect 7608 42950 7660 43002
rect 7672 42950 7724 43002
rect 7736 42950 7788 43002
rect 7800 42950 7852 43002
rect 7864 42950 7916 43002
rect 12047 42950 12099 43002
rect 12111 42950 12163 43002
rect 12175 42950 12227 43002
rect 12239 42950 12291 43002
rect 12303 42950 12355 43002
rect 16486 42950 16538 43002
rect 16550 42950 16602 43002
rect 16614 42950 16666 43002
rect 16678 42950 16730 43002
rect 16742 42950 16794 43002
rect 5388 42406 5440 42458
rect 5452 42406 5504 42458
rect 5516 42406 5568 42458
rect 5580 42406 5632 42458
rect 5644 42406 5696 42458
rect 9827 42406 9879 42458
rect 9891 42406 9943 42458
rect 9955 42406 10007 42458
rect 10019 42406 10071 42458
rect 10083 42406 10135 42458
rect 14266 42406 14318 42458
rect 14330 42406 14382 42458
rect 14394 42406 14446 42458
rect 14458 42406 14510 42458
rect 14522 42406 14574 42458
rect 18705 42406 18757 42458
rect 18769 42406 18821 42458
rect 18833 42406 18885 42458
rect 18897 42406 18949 42458
rect 18961 42406 19013 42458
rect 3169 41862 3221 41914
rect 3233 41862 3285 41914
rect 3297 41862 3349 41914
rect 3361 41862 3413 41914
rect 3425 41862 3477 41914
rect 7608 41862 7660 41914
rect 7672 41862 7724 41914
rect 7736 41862 7788 41914
rect 7800 41862 7852 41914
rect 7864 41862 7916 41914
rect 12047 41862 12099 41914
rect 12111 41862 12163 41914
rect 12175 41862 12227 41914
rect 12239 41862 12291 41914
rect 12303 41862 12355 41914
rect 16486 41862 16538 41914
rect 16550 41862 16602 41914
rect 16614 41862 16666 41914
rect 16678 41862 16730 41914
rect 16742 41862 16794 41914
rect 5388 41318 5440 41370
rect 5452 41318 5504 41370
rect 5516 41318 5568 41370
rect 5580 41318 5632 41370
rect 5644 41318 5696 41370
rect 9827 41318 9879 41370
rect 9891 41318 9943 41370
rect 9955 41318 10007 41370
rect 10019 41318 10071 41370
rect 10083 41318 10135 41370
rect 14266 41318 14318 41370
rect 14330 41318 14382 41370
rect 14394 41318 14446 41370
rect 14458 41318 14510 41370
rect 14522 41318 14574 41370
rect 18705 41318 18757 41370
rect 18769 41318 18821 41370
rect 18833 41318 18885 41370
rect 18897 41318 18949 41370
rect 18961 41318 19013 41370
rect 2504 41080 2556 41132
rect 940 40944 992 40996
rect 3169 40774 3221 40826
rect 3233 40774 3285 40826
rect 3297 40774 3349 40826
rect 3361 40774 3413 40826
rect 3425 40774 3477 40826
rect 7608 40774 7660 40826
rect 7672 40774 7724 40826
rect 7736 40774 7788 40826
rect 7800 40774 7852 40826
rect 7864 40774 7916 40826
rect 12047 40774 12099 40826
rect 12111 40774 12163 40826
rect 12175 40774 12227 40826
rect 12239 40774 12291 40826
rect 12303 40774 12355 40826
rect 16486 40774 16538 40826
rect 16550 40774 16602 40826
rect 16614 40774 16666 40826
rect 16678 40774 16730 40826
rect 16742 40774 16794 40826
rect 5388 40230 5440 40282
rect 5452 40230 5504 40282
rect 5516 40230 5568 40282
rect 5580 40230 5632 40282
rect 5644 40230 5696 40282
rect 9827 40230 9879 40282
rect 9891 40230 9943 40282
rect 9955 40230 10007 40282
rect 10019 40230 10071 40282
rect 10083 40230 10135 40282
rect 14266 40230 14318 40282
rect 14330 40230 14382 40282
rect 14394 40230 14446 40282
rect 14458 40230 14510 40282
rect 14522 40230 14574 40282
rect 18705 40230 18757 40282
rect 18769 40230 18821 40282
rect 18833 40230 18885 40282
rect 18897 40230 18949 40282
rect 18961 40230 19013 40282
rect 3169 39686 3221 39738
rect 3233 39686 3285 39738
rect 3297 39686 3349 39738
rect 3361 39686 3413 39738
rect 3425 39686 3477 39738
rect 7608 39686 7660 39738
rect 7672 39686 7724 39738
rect 7736 39686 7788 39738
rect 7800 39686 7852 39738
rect 7864 39686 7916 39738
rect 12047 39686 12099 39738
rect 12111 39686 12163 39738
rect 12175 39686 12227 39738
rect 12239 39686 12291 39738
rect 12303 39686 12355 39738
rect 16486 39686 16538 39738
rect 16550 39686 16602 39738
rect 16614 39686 16666 39738
rect 16678 39686 16730 39738
rect 16742 39686 16794 39738
rect 5388 39142 5440 39194
rect 5452 39142 5504 39194
rect 5516 39142 5568 39194
rect 5580 39142 5632 39194
rect 5644 39142 5696 39194
rect 9827 39142 9879 39194
rect 9891 39142 9943 39194
rect 9955 39142 10007 39194
rect 10019 39142 10071 39194
rect 10083 39142 10135 39194
rect 14266 39142 14318 39194
rect 14330 39142 14382 39194
rect 14394 39142 14446 39194
rect 14458 39142 14510 39194
rect 14522 39142 14574 39194
rect 18705 39142 18757 39194
rect 18769 39142 18821 39194
rect 18833 39142 18885 39194
rect 18897 39142 18949 39194
rect 18961 39142 19013 39194
rect 3169 38598 3221 38650
rect 3233 38598 3285 38650
rect 3297 38598 3349 38650
rect 3361 38598 3413 38650
rect 3425 38598 3477 38650
rect 7608 38598 7660 38650
rect 7672 38598 7724 38650
rect 7736 38598 7788 38650
rect 7800 38598 7852 38650
rect 7864 38598 7916 38650
rect 12047 38598 12099 38650
rect 12111 38598 12163 38650
rect 12175 38598 12227 38650
rect 12239 38598 12291 38650
rect 12303 38598 12355 38650
rect 16486 38598 16538 38650
rect 16550 38598 16602 38650
rect 16614 38598 16666 38650
rect 16678 38598 16730 38650
rect 16742 38598 16794 38650
rect 5388 38054 5440 38106
rect 5452 38054 5504 38106
rect 5516 38054 5568 38106
rect 5580 38054 5632 38106
rect 5644 38054 5696 38106
rect 9827 38054 9879 38106
rect 9891 38054 9943 38106
rect 9955 38054 10007 38106
rect 10019 38054 10071 38106
rect 10083 38054 10135 38106
rect 14266 38054 14318 38106
rect 14330 38054 14382 38106
rect 14394 38054 14446 38106
rect 14458 38054 14510 38106
rect 14522 38054 14574 38106
rect 18705 38054 18757 38106
rect 18769 38054 18821 38106
rect 18833 38054 18885 38106
rect 18897 38054 18949 38106
rect 18961 38054 19013 38106
rect 940 37612 992 37664
rect 3169 37510 3221 37562
rect 3233 37510 3285 37562
rect 3297 37510 3349 37562
rect 3361 37510 3413 37562
rect 3425 37510 3477 37562
rect 7608 37510 7660 37562
rect 7672 37510 7724 37562
rect 7736 37510 7788 37562
rect 7800 37510 7852 37562
rect 7864 37510 7916 37562
rect 12047 37510 12099 37562
rect 12111 37510 12163 37562
rect 12175 37510 12227 37562
rect 12239 37510 12291 37562
rect 12303 37510 12355 37562
rect 16486 37510 16538 37562
rect 16550 37510 16602 37562
rect 16614 37510 16666 37562
rect 16678 37510 16730 37562
rect 16742 37510 16794 37562
rect 5388 36966 5440 37018
rect 5452 36966 5504 37018
rect 5516 36966 5568 37018
rect 5580 36966 5632 37018
rect 5644 36966 5696 37018
rect 9827 36966 9879 37018
rect 9891 36966 9943 37018
rect 9955 36966 10007 37018
rect 10019 36966 10071 37018
rect 10083 36966 10135 37018
rect 14266 36966 14318 37018
rect 14330 36966 14382 37018
rect 14394 36966 14446 37018
rect 14458 36966 14510 37018
rect 14522 36966 14574 37018
rect 18705 36966 18757 37018
rect 18769 36966 18821 37018
rect 18833 36966 18885 37018
rect 18897 36966 18949 37018
rect 18961 36966 19013 37018
rect 3169 36422 3221 36474
rect 3233 36422 3285 36474
rect 3297 36422 3349 36474
rect 3361 36422 3413 36474
rect 3425 36422 3477 36474
rect 7608 36422 7660 36474
rect 7672 36422 7724 36474
rect 7736 36422 7788 36474
rect 7800 36422 7852 36474
rect 7864 36422 7916 36474
rect 12047 36422 12099 36474
rect 12111 36422 12163 36474
rect 12175 36422 12227 36474
rect 12239 36422 12291 36474
rect 12303 36422 12355 36474
rect 16486 36422 16538 36474
rect 16550 36422 16602 36474
rect 16614 36422 16666 36474
rect 16678 36422 16730 36474
rect 16742 36422 16794 36474
rect 7288 36184 7340 36236
rect 4620 36048 4672 36100
rect 7196 36116 7248 36168
rect 6920 36048 6972 36100
rect 5388 35878 5440 35930
rect 5452 35878 5504 35930
rect 5516 35878 5568 35930
rect 5580 35878 5632 35930
rect 5644 35878 5696 35930
rect 9827 35878 9879 35930
rect 9891 35878 9943 35930
rect 9955 35878 10007 35930
rect 10019 35878 10071 35930
rect 10083 35878 10135 35930
rect 14266 35878 14318 35930
rect 14330 35878 14382 35930
rect 14394 35878 14446 35930
rect 14458 35878 14510 35930
rect 14522 35878 14574 35930
rect 18705 35878 18757 35930
rect 18769 35878 18821 35930
rect 18833 35878 18885 35930
rect 18897 35878 18949 35930
rect 18961 35878 19013 35930
rect 4620 35683 4672 35692
rect 4620 35649 4629 35683
rect 4629 35649 4663 35683
rect 4663 35649 4672 35683
rect 4620 35640 4672 35649
rect 6184 35640 6236 35692
rect 5264 35436 5316 35488
rect 3169 35334 3221 35386
rect 3233 35334 3285 35386
rect 3297 35334 3349 35386
rect 3361 35334 3413 35386
rect 3425 35334 3477 35386
rect 7608 35334 7660 35386
rect 7672 35334 7724 35386
rect 7736 35334 7788 35386
rect 7800 35334 7852 35386
rect 7864 35334 7916 35386
rect 12047 35334 12099 35386
rect 12111 35334 12163 35386
rect 12175 35334 12227 35386
rect 12239 35334 12291 35386
rect 12303 35334 12355 35386
rect 16486 35334 16538 35386
rect 16550 35334 16602 35386
rect 16614 35334 16666 35386
rect 16678 35334 16730 35386
rect 16742 35334 16794 35386
rect 6092 35071 6144 35080
rect 6092 35037 6101 35071
rect 6101 35037 6135 35071
rect 6135 35037 6144 35071
rect 6092 35028 6144 35037
rect 6920 35071 6972 35080
rect 6920 35037 6929 35071
rect 6929 35037 6963 35071
rect 6963 35037 6972 35071
rect 6920 35028 6972 35037
rect 6368 34935 6420 34944
rect 6368 34901 6377 34935
rect 6377 34901 6411 34935
rect 6411 34901 6420 34935
rect 6368 34892 6420 34901
rect 5388 34790 5440 34842
rect 5452 34790 5504 34842
rect 5516 34790 5568 34842
rect 5580 34790 5632 34842
rect 5644 34790 5696 34842
rect 9827 34790 9879 34842
rect 9891 34790 9943 34842
rect 9955 34790 10007 34842
rect 10019 34790 10071 34842
rect 10083 34790 10135 34842
rect 14266 34790 14318 34842
rect 14330 34790 14382 34842
rect 14394 34790 14446 34842
rect 14458 34790 14510 34842
rect 14522 34790 14574 34842
rect 18705 34790 18757 34842
rect 18769 34790 18821 34842
rect 18833 34790 18885 34842
rect 18897 34790 18949 34842
rect 18961 34790 19013 34842
rect 6920 34620 6972 34672
rect 6460 34552 6512 34604
rect 7288 34595 7340 34604
rect 7288 34561 7297 34595
rect 7297 34561 7331 34595
rect 7331 34561 7340 34595
rect 7288 34552 7340 34561
rect 6184 34348 6236 34400
rect 3169 34246 3221 34298
rect 3233 34246 3285 34298
rect 3297 34246 3349 34298
rect 3361 34246 3413 34298
rect 3425 34246 3477 34298
rect 7608 34246 7660 34298
rect 7672 34246 7724 34298
rect 7736 34246 7788 34298
rect 7800 34246 7852 34298
rect 7864 34246 7916 34298
rect 12047 34246 12099 34298
rect 12111 34246 12163 34298
rect 12175 34246 12227 34298
rect 12239 34246 12291 34298
rect 12303 34246 12355 34298
rect 16486 34246 16538 34298
rect 16550 34246 16602 34298
rect 16614 34246 16666 34298
rect 16678 34246 16730 34298
rect 16742 34246 16794 34298
rect 6368 34144 6420 34196
rect 7380 34144 7432 34196
rect 8668 34076 8720 34128
rect 5724 34008 5776 34060
rect 6184 34051 6236 34060
rect 6184 34017 6193 34051
rect 6193 34017 6227 34051
rect 6227 34017 6236 34051
rect 6184 34008 6236 34017
rect 7196 34008 7248 34060
rect 6460 33940 6512 33992
rect 7288 33940 7340 33992
rect 940 33872 992 33924
rect 1676 33872 1728 33924
rect 5388 33702 5440 33754
rect 5452 33702 5504 33754
rect 5516 33702 5568 33754
rect 5580 33702 5632 33754
rect 5644 33702 5696 33754
rect 9827 33702 9879 33754
rect 9891 33702 9943 33754
rect 9955 33702 10007 33754
rect 10019 33702 10071 33754
rect 10083 33702 10135 33754
rect 14266 33702 14318 33754
rect 14330 33702 14382 33754
rect 14394 33702 14446 33754
rect 14458 33702 14510 33754
rect 14522 33702 14574 33754
rect 18705 33702 18757 33754
rect 18769 33702 18821 33754
rect 18833 33702 18885 33754
rect 18897 33702 18949 33754
rect 18961 33702 19013 33754
rect 3169 33158 3221 33210
rect 3233 33158 3285 33210
rect 3297 33158 3349 33210
rect 3361 33158 3413 33210
rect 3425 33158 3477 33210
rect 7608 33158 7660 33210
rect 7672 33158 7724 33210
rect 7736 33158 7788 33210
rect 7800 33158 7852 33210
rect 7864 33158 7916 33210
rect 12047 33158 12099 33210
rect 12111 33158 12163 33210
rect 12175 33158 12227 33210
rect 12239 33158 12291 33210
rect 12303 33158 12355 33210
rect 16486 33158 16538 33210
rect 16550 33158 16602 33210
rect 16614 33158 16666 33210
rect 16678 33158 16730 33210
rect 16742 33158 16794 33210
rect 7196 33056 7248 33108
rect 6092 32988 6144 33040
rect 6184 32988 6236 33040
rect 6184 32852 6236 32904
rect 7104 32852 7156 32904
rect 7932 32759 7984 32768
rect 7932 32725 7941 32759
rect 7941 32725 7975 32759
rect 7975 32725 7984 32759
rect 7932 32716 7984 32725
rect 5388 32614 5440 32666
rect 5452 32614 5504 32666
rect 5516 32614 5568 32666
rect 5580 32614 5632 32666
rect 5644 32614 5696 32666
rect 9827 32614 9879 32666
rect 9891 32614 9943 32666
rect 9955 32614 10007 32666
rect 10019 32614 10071 32666
rect 10083 32614 10135 32666
rect 14266 32614 14318 32666
rect 14330 32614 14382 32666
rect 14394 32614 14446 32666
rect 14458 32614 14510 32666
rect 14522 32614 14574 32666
rect 18705 32614 18757 32666
rect 18769 32614 18821 32666
rect 18833 32614 18885 32666
rect 18897 32614 18949 32666
rect 18961 32614 19013 32666
rect 4620 32376 4672 32428
rect 5172 32419 5224 32428
rect 5172 32385 5181 32419
rect 5181 32385 5215 32419
rect 5215 32385 5224 32419
rect 5172 32376 5224 32385
rect 5724 32444 5776 32496
rect 6828 32376 6880 32428
rect 6920 32376 6972 32428
rect 6092 32240 6144 32292
rect 6644 32172 6696 32224
rect 3169 32070 3221 32122
rect 3233 32070 3285 32122
rect 3297 32070 3349 32122
rect 3361 32070 3413 32122
rect 3425 32070 3477 32122
rect 7608 32070 7660 32122
rect 7672 32070 7724 32122
rect 7736 32070 7788 32122
rect 7800 32070 7852 32122
rect 7864 32070 7916 32122
rect 12047 32070 12099 32122
rect 12111 32070 12163 32122
rect 12175 32070 12227 32122
rect 12239 32070 12291 32122
rect 12303 32070 12355 32122
rect 16486 32070 16538 32122
rect 16550 32070 16602 32122
rect 16614 32070 16666 32122
rect 16678 32070 16730 32122
rect 16742 32070 16794 32122
rect 5264 31807 5316 31816
rect 5264 31773 5273 31807
rect 5273 31773 5307 31807
rect 5307 31773 5316 31807
rect 5264 31764 5316 31773
rect 5908 31807 5960 31816
rect 5908 31773 5917 31807
rect 5917 31773 5951 31807
rect 5951 31773 5960 31807
rect 5908 31764 5960 31773
rect 4712 31696 4764 31748
rect 5388 31526 5440 31578
rect 5452 31526 5504 31578
rect 5516 31526 5568 31578
rect 5580 31526 5632 31578
rect 5644 31526 5696 31578
rect 9827 31526 9879 31578
rect 9891 31526 9943 31578
rect 9955 31526 10007 31578
rect 10019 31526 10071 31578
rect 10083 31526 10135 31578
rect 14266 31526 14318 31578
rect 14330 31526 14382 31578
rect 14394 31526 14446 31578
rect 14458 31526 14510 31578
rect 14522 31526 14574 31578
rect 18705 31526 18757 31578
rect 18769 31526 18821 31578
rect 18833 31526 18885 31578
rect 18897 31526 18949 31578
rect 18961 31526 19013 31578
rect 5908 31467 5960 31476
rect 5908 31433 5917 31467
rect 5917 31433 5951 31467
rect 5951 31433 5960 31467
rect 5908 31424 5960 31433
rect 6460 31356 6512 31408
rect 5632 31288 5684 31340
rect 6000 31331 6052 31340
rect 6000 31297 6009 31331
rect 6009 31297 6043 31331
rect 6043 31297 6052 31331
rect 6000 31288 6052 31297
rect 6368 31288 6420 31340
rect 6828 31331 6880 31340
rect 6828 31297 6837 31331
rect 6837 31297 6871 31331
rect 6871 31297 6880 31331
rect 6828 31288 6880 31297
rect 5172 31220 5224 31272
rect 7104 31331 7156 31340
rect 7104 31297 7113 31331
rect 7113 31297 7147 31331
rect 7147 31297 7156 31331
rect 7104 31288 7156 31297
rect 7288 31220 7340 31272
rect 8852 31084 8904 31136
rect 3169 30982 3221 31034
rect 3233 30982 3285 31034
rect 3297 30982 3349 31034
rect 3361 30982 3413 31034
rect 3425 30982 3477 31034
rect 7608 30982 7660 31034
rect 7672 30982 7724 31034
rect 7736 30982 7788 31034
rect 7800 30982 7852 31034
rect 7864 30982 7916 31034
rect 12047 30982 12099 31034
rect 12111 30982 12163 31034
rect 12175 30982 12227 31034
rect 12239 30982 12291 31034
rect 12303 30982 12355 31034
rect 16486 30982 16538 31034
rect 16550 30982 16602 31034
rect 16614 30982 16666 31034
rect 16678 30982 16730 31034
rect 16742 30982 16794 31034
rect 6460 30812 6512 30864
rect 5724 30744 5776 30796
rect 940 30676 992 30728
rect 6000 30719 6052 30728
rect 6000 30685 6009 30719
rect 6009 30685 6043 30719
rect 6043 30685 6052 30719
rect 6000 30676 6052 30685
rect 6368 30676 6420 30728
rect 6552 30608 6604 30660
rect 7196 30608 7248 30660
rect 7472 30719 7524 30728
rect 7472 30685 7481 30719
rect 7481 30685 7515 30719
rect 7515 30685 7524 30719
rect 7472 30676 7524 30685
rect 7564 30608 7616 30660
rect 6000 30540 6052 30592
rect 6920 30540 6972 30592
rect 8024 30540 8076 30592
rect 5388 30438 5440 30490
rect 5452 30438 5504 30490
rect 5516 30438 5568 30490
rect 5580 30438 5632 30490
rect 5644 30438 5696 30490
rect 9827 30438 9879 30490
rect 9891 30438 9943 30490
rect 9955 30438 10007 30490
rect 10019 30438 10071 30490
rect 10083 30438 10135 30490
rect 14266 30438 14318 30490
rect 14330 30438 14382 30490
rect 14394 30438 14446 30490
rect 14458 30438 14510 30490
rect 14522 30438 14574 30490
rect 18705 30438 18757 30490
rect 18769 30438 18821 30490
rect 18833 30438 18885 30490
rect 18897 30438 18949 30490
rect 18961 30438 19013 30490
rect 6736 30336 6788 30388
rect 7564 30336 7616 30388
rect 8944 30336 8996 30388
rect 6184 30268 6236 30320
rect 7012 30243 7064 30252
rect 7012 30209 7021 30243
rect 7021 30209 7055 30243
rect 7055 30209 7064 30243
rect 7012 30200 7064 30209
rect 7196 30132 7248 30184
rect 7932 30200 7984 30252
rect 7380 30107 7432 30116
rect 7380 30073 7389 30107
rect 7389 30073 7423 30107
rect 7423 30073 7432 30107
rect 7380 30064 7432 30073
rect 6828 29996 6880 30048
rect 8116 30039 8168 30048
rect 8116 30005 8125 30039
rect 8125 30005 8159 30039
rect 8159 30005 8168 30039
rect 8116 29996 8168 30005
rect 3169 29894 3221 29946
rect 3233 29894 3285 29946
rect 3297 29894 3349 29946
rect 3361 29894 3413 29946
rect 3425 29894 3477 29946
rect 7608 29894 7660 29946
rect 7672 29894 7724 29946
rect 7736 29894 7788 29946
rect 7800 29894 7852 29946
rect 7864 29894 7916 29946
rect 12047 29894 12099 29946
rect 12111 29894 12163 29946
rect 12175 29894 12227 29946
rect 12239 29894 12291 29946
rect 12303 29894 12355 29946
rect 16486 29894 16538 29946
rect 16550 29894 16602 29946
rect 16614 29894 16666 29946
rect 16678 29894 16730 29946
rect 16742 29894 16794 29946
rect 5724 29792 5776 29844
rect 7472 29835 7524 29844
rect 7472 29801 7481 29835
rect 7481 29801 7515 29835
rect 7515 29801 7524 29835
rect 7472 29792 7524 29801
rect 7012 29724 7064 29776
rect 8208 29724 8260 29776
rect 4988 29588 5040 29640
rect 6184 29631 6236 29640
rect 6184 29597 6193 29631
rect 6193 29597 6227 29631
rect 6227 29597 6236 29631
rect 6184 29588 6236 29597
rect 6736 29631 6788 29640
rect 6736 29597 6745 29631
rect 6745 29597 6779 29631
rect 6779 29597 6788 29631
rect 6736 29588 6788 29597
rect 7012 29588 7064 29640
rect 7380 29588 7432 29640
rect 5080 29520 5132 29572
rect 4620 29495 4672 29504
rect 4620 29461 4629 29495
rect 4629 29461 4663 29495
rect 4663 29461 4672 29495
rect 4620 29452 4672 29461
rect 4804 29495 4856 29504
rect 4804 29461 4813 29495
rect 4813 29461 4847 29495
rect 4847 29461 4856 29495
rect 4804 29452 4856 29461
rect 4896 29452 4948 29504
rect 5388 29350 5440 29402
rect 5452 29350 5504 29402
rect 5516 29350 5568 29402
rect 5580 29350 5632 29402
rect 5644 29350 5696 29402
rect 9827 29350 9879 29402
rect 9891 29350 9943 29402
rect 9955 29350 10007 29402
rect 10019 29350 10071 29402
rect 10083 29350 10135 29402
rect 14266 29350 14318 29402
rect 14330 29350 14382 29402
rect 14394 29350 14446 29402
rect 14458 29350 14510 29402
rect 14522 29350 14574 29402
rect 18705 29350 18757 29402
rect 18769 29350 18821 29402
rect 18833 29350 18885 29402
rect 18897 29350 18949 29402
rect 18961 29350 19013 29402
rect 6920 29248 6972 29300
rect 7472 29248 7524 29300
rect 4896 29180 4948 29232
rect 4528 29112 4580 29164
rect 4804 29044 4856 29096
rect 4988 29087 5040 29096
rect 4988 29053 4997 29087
rect 4997 29053 5031 29087
rect 5031 29053 5040 29087
rect 4988 29044 5040 29053
rect 5080 29087 5132 29096
rect 5080 29053 5089 29087
rect 5089 29053 5123 29087
rect 5123 29053 5132 29087
rect 5080 29044 5132 29053
rect 6644 29155 6696 29164
rect 6644 29121 6653 29155
rect 6653 29121 6687 29155
rect 6687 29121 6696 29155
rect 6644 29112 6696 29121
rect 6828 29155 6880 29164
rect 6828 29121 6837 29155
rect 6837 29121 6871 29155
rect 6871 29121 6880 29155
rect 6828 29112 6880 29121
rect 7104 29112 7156 29164
rect 7472 29112 7524 29164
rect 8024 29155 8076 29164
rect 8024 29121 8033 29155
rect 8033 29121 8067 29155
rect 8067 29121 8076 29155
rect 8024 29112 8076 29121
rect 6736 29044 6788 29096
rect 6460 28976 6512 29028
rect 4712 28951 4764 28960
rect 4712 28917 4721 28951
rect 4721 28917 4755 28951
rect 4755 28917 4764 28951
rect 4712 28908 4764 28917
rect 5264 28908 5316 28960
rect 3169 28806 3221 28858
rect 3233 28806 3285 28858
rect 3297 28806 3349 28858
rect 3361 28806 3413 28858
rect 3425 28806 3477 28858
rect 7608 28806 7660 28858
rect 7672 28806 7724 28858
rect 7736 28806 7788 28858
rect 7800 28806 7852 28858
rect 7864 28806 7916 28858
rect 12047 28806 12099 28858
rect 12111 28806 12163 28858
rect 12175 28806 12227 28858
rect 12239 28806 12291 28858
rect 12303 28806 12355 28858
rect 16486 28806 16538 28858
rect 16550 28806 16602 28858
rect 16614 28806 16666 28858
rect 16678 28806 16730 28858
rect 16742 28806 16794 28858
rect 4160 28704 4212 28756
rect 4620 28636 4672 28688
rect 5724 28636 5776 28688
rect 6460 28611 6512 28620
rect 6460 28577 6469 28611
rect 6469 28577 6503 28611
rect 6503 28577 6512 28611
rect 6460 28568 6512 28577
rect 6828 28568 6880 28620
rect 4068 28500 4120 28552
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6595 28543
rect 6595 28509 6604 28543
rect 6552 28500 6604 28509
rect 6736 28543 6788 28552
rect 6736 28509 6745 28543
rect 6745 28509 6779 28543
rect 6779 28509 6788 28543
rect 6736 28500 6788 28509
rect 7288 28500 7340 28552
rect 7472 28543 7524 28552
rect 7472 28509 7481 28543
rect 7481 28509 7515 28543
rect 7515 28509 7524 28543
rect 7472 28500 7524 28509
rect 7932 28500 7984 28552
rect 3792 28432 3844 28484
rect 4712 28432 4764 28484
rect 3976 28364 4028 28416
rect 4252 28407 4304 28416
rect 4252 28373 4261 28407
rect 4261 28373 4295 28407
rect 4295 28373 4304 28407
rect 4252 28364 4304 28373
rect 6276 28407 6328 28416
rect 6276 28373 6285 28407
rect 6285 28373 6319 28407
rect 6319 28373 6328 28407
rect 6276 28364 6328 28373
rect 7288 28364 7340 28416
rect 5388 28262 5440 28314
rect 5452 28262 5504 28314
rect 5516 28262 5568 28314
rect 5580 28262 5632 28314
rect 5644 28262 5696 28314
rect 9827 28262 9879 28314
rect 9891 28262 9943 28314
rect 9955 28262 10007 28314
rect 10019 28262 10071 28314
rect 10083 28262 10135 28314
rect 14266 28262 14318 28314
rect 14330 28262 14382 28314
rect 14394 28262 14446 28314
rect 14458 28262 14510 28314
rect 14522 28262 14574 28314
rect 18705 28262 18757 28314
rect 18769 28262 18821 28314
rect 18833 28262 18885 28314
rect 18897 28262 18949 28314
rect 18961 28262 19013 28314
rect 6460 28024 6512 28076
rect 8944 28024 8996 28076
rect 8024 27956 8076 28008
rect 3169 27718 3221 27770
rect 3233 27718 3285 27770
rect 3297 27718 3349 27770
rect 3361 27718 3413 27770
rect 3425 27718 3477 27770
rect 7608 27718 7660 27770
rect 7672 27718 7724 27770
rect 7736 27718 7788 27770
rect 7800 27718 7852 27770
rect 7864 27718 7916 27770
rect 12047 27718 12099 27770
rect 12111 27718 12163 27770
rect 12175 27718 12227 27770
rect 12239 27718 12291 27770
rect 12303 27718 12355 27770
rect 16486 27718 16538 27770
rect 16550 27718 16602 27770
rect 16614 27718 16666 27770
rect 16678 27718 16730 27770
rect 16742 27718 16794 27770
rect 4252 27548 4304 27600
rect 3608 27480 3660 27532
rect 5816 27480 5868 27532
rect 3792 27412 3844 27464
rect 4068 27412 4120 27464
rect 4436 27455 4488 27464
rect 4436 27421 4445 27455
rect 4445 27421 4479 27455
rect 4479 27421 4488 27455
rect 4436 27412 4488 27421
rect 4620 27455 4672 27464
rect 4620 27421 4629 27455
rect 4629 27421 4663 27455
rect 4663 27421 4672 27455
rect 4620 27412 4672 27421
rect 6828 27344 6880 27396
rect 6644 27276 6696 27328
rect 5388 27174 5440 27226
rect 5452 27174 5504 27226
rect 5516 27174 5568 27226
rect 5580 27174 5632 27226
rect 5644 27174 5696 27226
rect 9827 27174 9879 27226
rect 9891 27174 9943 27226
rect 9955 27174 10007 27226
rect 10019 27174 10071 27226
rect 10083 27174 10135 27226
rect 14266 27174 14318 27226
rect 14330 27174 14382 27226
rect 14394 27174 14446 27226
rect 14458 27174 14510 27226
rect 14522 27174 14574 27226
rect 18705 27174 18757 27226
rect 18769 27174 18821 27226
rect 18833 27174 18885 27226
rect 18897 27174 18949 27226
rect 18961 27174 19013 27226
rect 3608 27072 3660 27124
rect 4160 27072 4212 27124
rect 4988 27072 5040 27124
rect 2872 27004 2924 27056
rect 4068 27004 4120 27056
rect 6184 27004 6236 27056
rect 6828 27004 6880 27056
rect 7472 27004 7524 27056
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 4344 26936 4396 26988
rect 5632 26979 5684 26988
rect 5632 26945 5641 26979
rect 5641 26945 5675 26979
rect 5675 26945 5684 26979
rect 5632 26936 5684 26945
rect 6368 26936 6420 26988
rect 2136 26868 2188 26920
rect 4896 26868 4948 26920
rect 6920 26868 6972 26920
rect 7380 26868 7432 26920
rect 940 26800 992 26852
rect 6736 26800 6788 26852
rect 8300 26843 8352 26852
rect 8300 26809 8309 26843
rect 8309 26809 8343 26843
rect 8343 26809 8352 26843
rect 8300 26800 8352 26809
rect 5908 26775 5960 26784
rect 5908 26741 5917 26775
rect 5917 26741 5951 26775
rect 5951 26741 5960 26775
rect 5908 26732 5960 26741
rect 8484 26775 8536 26784
rect 8484 26741 8493 26775
rect 8493 26741 8527 26775
rect 8527 26741 8536 26775
rect 8484 26732 8536 26741
rect 3169 26630 3221 26682
rect 3233 26630 3285 26682
rect 3297 26630 3349 26682
rect 3361 26630 3413 26682
rect 3425 26630 3477 26682
rect 7608 26630 7660 26682
rect 7672 26630 7724 26682
rect 7736 26630 7788 26682
rect 7800 26630 7852 26682
rect 7864 26630 7916 26682
rect 12047 26630 12099 26682
rect 12111 26630 12163 26682
rect 12175 26630 12227 26682
rect 12239 26630 12291 26682
rect 12303 26630 12355 26682
rect 16486 26630 16538 26682
rect 16550 26630 16602 26682
rect 16614 26630 16666 26682
rect 16678 26630 16730 26682
rect 16742 26630 16794 26682
rect 4436 26528 4488 26580
rect 4528 26571 4580 26580
rect 4528 26537 4537 26571
rect 4537 26537 4571 26571
rect 4571 26537 4580 26571
rect 4528 26528 4580 26537
rect 4712 26460 4764 26512
rect 6276 26460 6328 26512
rect 8760 26460 8812 26512
rect 2596 26392 2648 26444
rect 4344 26392 4396 26444
rect 6092 26392 6144 26444
rect 4896 26367 4948 26376
rect 4896 26333 4905 26367
rect 4905 26333 4939 26367
rect 4939 26333 4948 26367
rect 4896 26324 4948 26333
rect 5816 26367 5868 26376
rect 5816 26333 5825 26367
rect 5825 26333 5859 26367
rect 5859 26333 5868 26367
rect 5816 26324 5868 26333
rect 6000 26367 6052 26376
rect 6000 26333 6009 26367
rect 6009 26333 6043 26367
rect 6043 26333 6052 26367
rect 6000 26324 6052 26333
rect 6460 26324 6512 26376
rect 2044 26188 2096 26240
rect 5080 26256 5132 26308
rect 6184 26299 6236 26308
rect 6184 26265 6193 26299
rect 6193 26265 6227 26299
rect 6227 26265 6236 26299
rect 6184 26256 6236 26265
rect 7288 26324 7340 26376
rect 7932 26256 7984 26308
rect 8576 26256 8628 26308
rect 8208 26188 8260 26240
rect 8392 26188 8444 26240
rect 5388 26086 5440 26138
rect 5452 26086 5504 26138
rect 5516 26086 5568 26138
rect 5580 26086 5632 26138
rect 5644 26086 5696 26138
rect 9827 26086 9879 26138
rect 9891 26086 9943 26138
rect 9955 26086 10007 26138
rect 10019 26086 10071 26138
rect 10083 26086 10135 26138
rect 14266 26086 14318 26138
rect 14330 26086 14382 26138
rect 14394 26086 14446 26138
rect 14458 26086 14510 26138
rect 14522 26086 14574 26138
rect 18705 26086 18757 26138
rect 18769 26086 18821 26138
rect 18833 26086 18885 26138
rect 18897 26086 18949 26138
rect 18961 26086 19013 26138
rect 7012 25984 7064 26036
rect 4436 25916 4488 25968
rect 4344 25848 4396 25900
rect 4620 25848 4672 25900
rect 6828 25916 6880 25968
rect 5080 25780 5132 25832
rect 7472 25848 7524 25900
rect 6920 25823 6972 25832
rect 6920 25789 6929 25823
rect 6929 25789 6963 25823
rect 6963 25789 6972 25823
rect 6920 25780 6972 25789
rect 7380 25780 7432 25832
rect 5172 25644 5224 25696
rect 3169 25542 3221 25594
rect 3233 25542 3285 25594
rect 3297 25542 3349 25594
rect 3361 25542 3413 25594
rect 3425 25542 3477 25594
rect 7608 25542 7660 25594
rect 7672 25542 7724 25594
rect 7736 25542 7788 25594
rect 7800 25542 7852 25594
rect 7864 25542 7916 25594
rect 12047 25542 12099 25594
rect 12111 25542 12163 25594
rect 12175 25542 12227 25594
rect 12239 25542 12291 25594
rect 12303 25542 12355 25594
rect 16486 25542 16538 25594
rect 16550 25542 16602 25594
rect 16614 25542 16666 25594
rect 16678 25542 16730 25594
rect 16742 25542 16794 25594
rect 2136 25483 2188 25492
rect 2136 25449 2145 25483
rect 2145 25449 2179 25483
rect 2179 25449 2188 25483
rect 2136 25440 2188 25449
rect 5816 25440 5868 25492
rect 5724 25372 5776 25424
rect 8116 25483 8168 25492
rect 8116 25449 8125 25483
rect 8125 25449 8159 25483
rect 8159 25449 8168 25483
rect 8116 25440 8168 25449
rect 7012 25304 7064 25356
rect 3608 25236 3660 25288
rect 4068 25236 4120 25288
rect 5816 25279 5868 25288
rect 5816 25245 5825 25279
rect 5825 25245 5859 25279
rect 5859 25245 5868 25279
rect 5816 25236 5868 25245
rect 7840 25279 7892 25288
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 7840 25236 7892 25245
rect 2044 25168 2096 25220
rect 6368 25168 6420 25220
rect 6828 25168 6880 25220
rect 8300 25211 8352 25220
rect 8300 25177 8309 25211
rect 8309 25177 8343 25211
rect 8343 25177 8352 25211
rect 8300 25168 8352 25177
rect 1952 25143 2004 25152
rect 1952 25109 1961 25143
rect 1961 25109 1995 25143
rect 1995 25109 2004 25143
rect 1952 25100 2004 25109
rect 2228 25100 2280 25152
rect 6736 25100 6788 25152
rect 8208 25100 8260 25152
rect 5388 24998 5440 25050
rect 5452 24998 5504 25050
rect 5516 24998 5568 25050
rect 5580 24998 5632 25050
rect 5644 24998 5696 25050
rect 9827 24998 9879 25050
rect 9891 24998 9943 25050
rect 9955 24998 10007 25050
rect 10019 24998 10071 25050
rect 10083 24998 10135 25050
rect 14266 24998 14318 25050
rect 14330 24998 14382 25050
rect 14394 24998 14446 25050
rect 14458 24998 14510 25050
rect 14522 24998 14574 25050
rect 18705 24998 18757 25050
rect 18769 24998 18821 25050
rect 18833 24998 18885 25050
rect 18897 24998 18949 25050
rect 18961 24998 19013 25050
rect 4068 24896 4120 24948
rect 5080 24896 5132 24948
rect 6828 24828 6880 24880
rect 4896 24760 4948 24812
rect 2228 24692 2280 24744
rect 4804 24692 4856 24744
rect 6644 24692 6696 24744
rect 8392 24828 8444 24880
rect 9128 24828 9180 24880
rect 8024 24760 8076 24812
rect 7932 24692 7984 24744
rect 2688 24556 2740 24608
rect 7104 24624 7156 24676
rect 4160 24556 4212 24608
rect 7472 24556 7524 24608
rect 7564 24556 7616 24608
rect 3169 24454 3221 24506
rect 3233 24454 3285 24506
rect 3297 24454 3349 24506
rect 3361 24454 3413 24506
rect 3425 24454 3477 24506
rect 7608 24454 7660 24506
rect 7672 24454 7724 24506
rect 7736 24454 7788 24506
rect 7800 24454 7852 24506
rect 7864 24454 7916 24506
rect 12047 24454 12099 24506
rect 12111 24454 12163 24506
rect 12175 24454 12227 24506
rect 12239 24454 12291 24506
rect 12303 24454 12355 24506
rect 16486 24454 16538 24506
rect 16550 24454 16602 24506
rect 16614 24454 16666 24506
rect 16678 24454 16730 24506
rect 16742 24454 16794 24506
rect 4160 24395 4212 24404
rect 4160 24361 4169 24395
rect 4169 24361 4203 24395
rect 4203 24361 4212 24395
rect 4160 24352 4212 24361
rect 2228 24216 2280 24268
rect 2136 24191 2188 24200
rect 2136 24157 2145 24191
rect 2145 24157 2179 24191
rect 2179 24157 2188 24191
rect 2136 24148 2188 24157
rect 6276 24352 6328 24404
rect 6736 24352 6788 24404
rect 7840 24352 7892 24404
rect 5816 24284 5868 24336
rect 1032 24080 1084 24132
rect 4988 24148 5040 24200
rect 7012 24216 7064 24268
rect 6092 24148 6144 24200
rect 6552 24148 6604 24200
rect 7288 24148 7340 24200
rect 7840 24148 7892 24200
rect 5816 24080 5868 24132
rect 9680 24080 9732 24132
rect 2044 24012 2096 24064
rect 2964 24012 3016 24064
rect 4344 24012 4396 24064
rect 9036 24012 9088 24064
rect 5388 23910 5440 23962
rect 5452 23910 5504 23962
rect 5516 23910 5568 23962
rect 5580 23910 5632 23962
rect 5644 23910 5696 23962
rect 9827 23910 9879 23962
rect 9891 23910 9943 23962
rect 9955 23910 10007 23962
rect 10019 23910 10071 23962
rect 10083 23910 10135 23962
rect 14266 23910 14318 23962
rect 14330 23910 14382 23962
rect 14394 23910 14446 23962
rect 14458 23910 14510 23962
rect 14522 23910 14574 23962
rect 18705 23910 18757 23962
rect 18769 23910 18821 23962
rect 18833 23910 18885 23962
rect 18897 23910 18949 23962
rect 18961 23910 19013 23962
rect 4068 23808 4120 23860
rect 4344 23808 4396 23860
rect 4712 23808 4764 23860
rect 6368 23808 6420 23860
rect 4068 23715 4120 23724
rect 4068 23681 4077 23715
rect 4077 23681 4111 23715
rect 4111 23681 4120 23715
rect 4068 23672 4120 23681
rect 4252 23715 4304 23724
rect 4252 23681 4261 23715
rect 4261 23681 4295 23715
rect 4295 23681 4304 23715
rect 4252 23672 4304 23681
rect 4712 23672 4764 23724
rect 5264 23672 5316 23724
rect 7104 23715 7156 23724
rect 7104 23681 7113 23715
rect 7113 23681 7147 23715
rect 7147 23681 7156 23715
rect 7104 23672 7156 23681
rect 7472 23672 7524 23724
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 6552 23604 6604 23656
rect 4252 23536 4304 23588
rect 940 23468 992 23520
rect 3169 23366 3221 23418
rect 3233 23366 3285 23418
rect 3297 23366 3349 23418
rect 3361 23366 3413 23418
rect 3425 23366 3477 23418
rect 7608 23366 7660 23418
rect 7672 23366 7724 23418
rect 7736 23366 7788 23418
rect 7800 23366 7852 23418
rect 7864 23366 7916 23418
rect 12047 23366 12099 23418
rect 12111 23366 12163 23418
rect 12175 23366 12227 23418
rect 12239 23366 12291 23418
rect 12303 23366 12355 23418
rect 16486 23366 16538 23418
rect 16550 23366 16602 23418
rect 16614 23366 16666 23418
rect 16678 23366 16730 23418
rect 16742 23366 16794 23418
rect 5908 23307 5960 23316
rect 5908 23273 5917 23307
rect 5917 23273 5951 23307
rect 5951 23273 5960 23307
rect 5908 23264 5960 23273
rect 6000 23196 6052 23248
rect 6184 23128 6236 23180
rect 8300 23264 8352 23316
rect 6000 23103 6052 23112
rect 6000 23069 6009 23103
rect 6009 23069 6043 23103
rect 6043 23069 6052 23103
rect 6000 23060 6052 23069
rect 6552 23035 6604 23044
rect 6552 23001 6561 23035
rect 6561 23001 6595 23035
rect 6595 23001 6604 23035
rect 6552 22992 6604 23001
rect 7104 22924 7156 22976
rect 8300 22924 8352 22976
rect 5388 22822 5440 22874
rect 5452 22822 5504 22874
rect 5516 22822 5568 22874
rect 5580 22822 5632 22874
rect 5644 22822 5696 22874
rect 9827 22822 9879 22874
rect 9891 22822 9943 22874
rect 9955 22822 10007 22874
rect 10019 22822 10071 22874
rect 10083 22822 10135 22874
rect 14266 22822 14318 22874
rect 14330 22822 14382 22874
rect 14394 22822 14446 22874
rect 14458 22822 14510 22874
rect 14522 22822 14574 22874
rect 18705 22822 18757 22874
rect 18769 22822 18821 22874
rect 18833 22822 18885 22874
rect 18897 22822 18949 22874
rect 18961 22822 19013 22874
rect 5724 22763 5776 22772
rect 5724 22729 5733 22763
rect 5733 22729 5767 22763
rect 5767 22729 5776 22763
rect 5724 22720 5776 22729
rect 6000 22720 6052 22772
rect 6828 22720 6880 22772
rect 7288 22720 7340 22772
rect 8116 22720 8168 22772
rect 8300 22720 8352 22772
rect 1768 22652 1820 22704
rect 2596 22652 2648 22704
rect 4068 22652 4120 22704
rect 6368 22652 6420 22704
rect 7380 22652 7432 22704
rect 1952 22584 2004 22636
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 6644 22584 6696 22636
rect 7104 22627 7156 22636
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 7104 22584 7156 22593
rect 7472 22584 7524 22636
rect 1860 22559 1912 22568
rect 1860 22525 1869 22559
rect 1869 22525 1903 22559
rect 1903 22525 1912 22559
rect 1860 22516 1912 22525
rect 8300 22627 8352 22636
rect 8300 22593 8309 22627
rect 8309 22593 8343 22627
rect 8343 22593 8352 22627
rect 8300 22584 8352 22593
rect 8944 22584 8996 22636
rect 2136 22380 2188 22432
rect 7472 22380 7524 22432
rect 7840 22380 7892 22432
rect 7932 22380 7984 22432
rect 3169 22278 3221 22330
rect 3233 22278 3285 22330
rect 3297 22278 3349 22330
rect 3361 22278 3413 22330
rect 3425 22278 3477 22330
rect 7608 22278 7660 22330
rect 7672 22278 7724 22330
rect 7736 22278 7788 22330
rect 7800 22278 7852 22330
rect 7864 22278 7916 22330
rect 12047 22278 12099 22330
rect 12111 22278 12163 22330
rect 12175 22278 12227 22330
rect 12239 22278 12291 22330
rect 12303 22278 12355 22330
rect 16486 22278 16538 22330
rect 16550 22278 16602 22330
rect 16614 22278 16666 22330
rect 16678 22278 16730 22330
rect 16742 22278 16794 22330
rect 4436 22219 4488 22228
rect 4436 22185 4445 22219
rect 4445 22185 4479 22219
rect 4479 22185 4488 22219
rect 4436 22176 4488 22185
rect 5724 22176 5776 22228
rect 7104 22176 7156 22228
rect 7196 22176 7248 22228
rect 8116 22176 8168 22228
rect 1860 21904 1912 21956
rect 2780 21904 2832 21956
rect 6184 22040 6236 22092
rect 4988 21972 5040 22024
rect 6092 21972 6144 22024
rect 7104 21972 7156 22024
rect 4804 21904 4856 21956
rect 5724 21904 5776 21956
rect 5816 21947 5868 21956
rect 5816 21913 5825 21947
rect 5825 21913 5859 21947
rect 5859 21913 5868 21947
rect 5816 21904 5868 21913
rect 6184 21904 6236 21956
rect 7380 21904 7432 21956
rect 7840 21947 7892 21956
rect 7840 21913 7849 21947
rect 7849 21913 7883 21947
rect 7883 21913 7892 21947
rect 7840 21904 7892 21913
rect 8208 21904 8260 21956
rect 1584 21836 1636 21888
rect 5264 21836 5316 21888
rect 6092 21836 6144 21888
rect 6368 21836 6420 21888
rect 5388 21734 5440 21786
rect 5452 21734 5504 21786
rect 5516 21734 5568 21786
rect 5580 21734 5632 21786
rect 5644 21734 5696 21786
rect 9827 21734 9879 21786
rect 9891 21734 9943 21786
rect 9955 21734 10007 21786
rect 10019 21734 10071 21786
rect 10083 21734 10135 21786
rect 14266 21734 14318 21786
rect 14330 21734 14382 21786
rect 14394 21734 14446 21786
rect 14458 21734 14510 21786
rect 14522 21734 14574 21786
rect 18705 21734 18757 21786
rect 18769 21734 18821 21786
rect 18833 21734 18885 21786
rect 18897 21734 18949 21786
rect 18961 21734 19013 21786
rect 5264 21632 5316 21684
rect 6092 21632 6144 21684
rect 5908 21564 5960 21616
rect 4988 21496 5040 21548
rect 5264 21496 5316 21548
rect 5724 21539 5776 21548
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 7840 21564 7892 21616
rect 5908 21428 5960 21480
rect 8208 21496 8260 21548
rect 8944 21428 8996 21480
rect 8392 21360 8444 21412
rect 8300 21292 8352 21344
rect 3169 21190 3221 21242
rect 3233 21190 3285 21242
rect 3297 21190 3349 21242
rect 3361 21190 3413 21242
rect 3425 21190 3477 21242
rect 7608 21190 7660 21242
rect 7672 21190 7724 21242
rect 7736 21190 7788 21242
rect 7800 21190 7852 21242
rect 7864 21190 7916 21242
rect 12047 21190 12099 21242
rect 12111 21190 12163 21242
rect 12175 21190 12227 21242
rect 12239 21190 12291 21242
rect 12303 21190 12355 21242
rect 16486 21190 16538 21242
rect 16550 21190 16602 21242
rect 16614 21190 16666 21242
rect 16678 21190 16730 21242
rect 16742 21190 16794 21242
rect 2228 21088 2280 21140
rect 5080 21131 5132 21140
rect 5080 21097 5089 21131
rect 5089 21097 5123 21131
rect 5123 21097 5132 21131
rect 5080 21088 5132 21097
rect 8208 21131 8260 21140
rect 8208 21097 8217 21131
rect 8217 21097 8251 21131
rect 8251 21097 8260 21131
rect 8208 21088 8260 21097
rect 2780 20952 2832 21004
rect 2044 20884 2096 20936
rect 2228 20884 2280 20936
rect 3700 20884 3752 20936
rect 5172 20884 5224 20936
rect 7472 20884 7524 20936
rect 3056 20816 3108 20868
rect 3976 20816 4028 20868
rect 5908 20816 5960 20868
rect 1860 20791 1912 20800
rect 1860 20757 1869 20791
rect 1869 20757 1903 20791
rect 1903 20757 1912 20791
rect 1860 20748 1912 20757
rect 3148 20791 3200 20800
rect 3148 20757 3157 20791
rect 3157 20757 3191 20791
rect 3191 20757 3200 20791
rect 3148 20748 3200 20757
rect 7196 20748 7248 20800
rect 7472 20748 7524 20800
rect 5388 20646 5440 20698
rect 5452 20646 5504 20698
rect 5516 20646 5568 20698
rect 5580 20646 5632 20698
rect 5644 20646 5696 20698
rect 9827 20646 9879 20698
rect 9891 20646 9943 20698
rect 9955 20646 10007 20698
rect 10019 20646 10071 20698
rect 10083 20646 10135 20698
rect 14266 20646 14318 20698
rect 14330 20646 14382 20698
rect 14394 20646 14446 20698
rect 14458 20646 14510 20698
rect 14522 20646 14574 20698
rect 18705 20646 18757 20698
rect 18769 20646 18821 20698
rect 18833 20646 18885 20698
rect 18897 20646 18949 20698
rect 18961 20646 19013 20698
rect 4436 20544 4488 20596
rect 5724 20476 5776 20528
rect 6092 20476 6144 20528
rect 3148 20408 3200 20460
rect 5264 20451 5316 20460
rect 5264 20417 5273 20451
rect 5273 20417 5307 20451
rect 5307 20417 5316 20451
rect 5264 20408 5316 20417
rect 5816 20408 5868 20460
rect 6368 20408 6420 20460
rect 3056 20340 3108 20392
rect 6276 20340 6328 20392
rect 6552 20340 6604 20392
rect 3700 20204 3752 20256
rect 6552 20204 6604 20256
rect 3169 20102 3221 20154
rect 3233 20102 3285 20154
rect 3297 20102 3349 20154
rect 3361 20102 3413 20154
rect 3425 20102 3477 20154
rect 7608 20102 7660 20154
rect 7672 20102 7724 20154
rect 7736 20102 7788 20154
rect 7800 20102 7852 20154
rect 7864 20102 7916 20154
rect 12047 20102 12099 20154
rect 12111 20102 12163 20154
rect 12175 20102 12227 20154
rect 12239 20102 12291 20154
rect 12303 20102 12355 20154
rect 16486 20102 16538 20154
rect 16550 20102 16602 20154
rect 16614 20102 16666 20154
rect 16678 20102 16730 20154
rect 16742 20102 16794 20154
rect 2964 20043 3016 20052
rect 2964 20009 2973 20043
rect 2973 20009 3007 20043
rect 3007 20009 3016 20043
rect 2964 20000 3016 20009
rect 1952 19932 2004 19984
rect 1216 19796 1268 19848
rect 940 19728 992 19780
rect 2780 19728 2832 19780
rect 3976 19728 4028 19780
rect 4068 19660 4120 19712
rect 5388 19558 5440 19610
rect 5452 19558 5504 19610
rect 5516 19558 5568 19610
rect 5580 19558 5632 19610
rect 5644 19558 5696 19610
rect 9827 19558 9879 19610
rect 9891 19558 9943 19610
rect 9955 19558 10007 19610
rect 10019 19558 10071 19610
rect 10083 19558 10135 19610
rect 14266 19558 14318 19610
rect 14330 19558 14382 19610
rect 14394 19558 14446 19610
rect 14458 19558 14510 19610
rect 14522 19558 14574 19610
rect 18705 19558 18757 19610
rect 18769 19558 18821 19610
rect 18833 19558 18885 19610
rect 18897 19558 18949 19610
rect 18961 19558 19013 19610
rect 4436 19456 4488 19508
rect 1860 19388 1912 19440
rect 1492 19320 1544 19372
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 2044 19320 2096 19329
rect 2136 19363 2188 19372
rect 2136 19329 2145 19363
rect 2145 19329 2179 19363
rect 2179 19329 2188 19363
rect 2136 19320 2188 19329
rect 2228 19320 2280 19372
rect 5724 19388 5776 19440
rect 4804 19320 4856 19372
rect 1952 19252 2004 19304
rect 3169 19014 3221 19066
rect 3233 19014 3285 19066
rect 3297 19014 3349 19066
rect 3361 19014 3413 19066
rect 3425 19014 3477 19066
rect 7608 19014 7660 19066
rect 7672 19014 7724 19066
rect 7736 19014 7788 19066
rect 7800 19014 7852 19066
rect 7864 19014 7916 19066
rect 12047 19014 12099 19066
rect 12111 19014 12163 19066
rect 12175 19014 12227 19066
rect 12239 19014 12291 19066
rect 12303 19014 12355 19066
rect 16486 19014 16538 19066
rect 16550 19014 16602 19066
rect 16614 19014 16666 19066
rect 16678 19014 16730 19066
rect 16742 19014 16794 19066
rect 3056 18912 3108 18964
rect 2780 18776 2832 18828
rect 3792 18912 3844 18964
rect 6460 18912 6512 18964
rect 2320 18708 2372 18760
rect 3240 18708 3292 18760
rect 3608 18640 3660 18692
rect 5908 18708 5960 18760
rect 6644 18640 6696 18692
rect 6920 18640 6972 18692
rect 5388 18470 5440 18522
rect 5452 18470 5504 18522
rect 5516 18470 5568 18522
rect 5580 18470 5632 18522
rect 5644 18470 5696 18522
rect 9827 18470 9879 18522
rect 9891 18470 9943 18522
rect 9955 18470 10007 18522
rect 10019 18470 10071 18522
rect 10083 18470 10135 18522
rect 14266 18470 14318 18522
rect 14330 18470 14382 18522
rect 14394 18470 14446 18522
rect 14458 18470 14510 18522
rect 14522 18470 14574 18522
rect 18705 18470 18757 18522
rect 18769 18470 18821 18522
rect 18833 18470 18885 18522
rect 18897 18470 18949 18522
rect 18961 18470 19013 18522
rect 2412 18232 2464 18284
rect 3240 18232 3292 18284
rect 4804 18232 4856 18284
rect 2320 18164 2372 18216
rect 2872 18096 2924 18148
rect 2504 18028 2556 18080
rect 3056 18028 3108 18080
rect 3169 17926 3221 17978
rect 3233 17926 3285 17978
rect 3297 17926 3349 17978
rect 3361 17926 3413 17978
rect 3425 17926 3477 17978
rect 7608 17926 7660 17978
rect 7672 17926 7724 17978
rect 7736 17926 7788 17978
rect 7800 17926 7852 17978
rect 7864 17926 7916 17978
rect 12047 17926 12099 17978
rect 12111 17926 12163 17978
rect 12175 17926 12227 17978
rect 12239 17926 12291 17978
rect 12303 17926 12355 17978
rect 16486 17926 16538 17978
rect 16550 17926 16602 17978
rect 16614 17926 16666 17978
rect 16678 17926 16730 17978
rect 16742 17926 16794 17978
rect 1860 17824 1912 17876
rect 2596 17824 2648 17876
rect 2964 17867 3016 17876
rect 2964 17833 2973 17867
rect 2973 17833 3007 17867
rect 3007 17833 3016 17867
rect 2964 17824 3016 17833
rect 3516 17824 3568 17876
rect 2228 17620 2280 17672
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 2136 17527 2188 17536
rect 2136 17493 2145 17527
rect 2145 17493 2179 17527
rect 2179 17493 2188 17527
rect 2136 17484 2188 17493
rect 2596 17484 2648 17536
rect 3884 17688 3936 17740
rect 3516 17620 3568 17672
rect 3700 17552 3752 17604
rect 3976 17484 4028 17536
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 5644 17382 5696 17434
rect 9827 17382 9879 17434
rect 9891 17382 9943 17434
rect 9955 17382 10007 17434
rect 10019 17382 10071 17434
rect 10083 17382 10135 17434
rect 14266 17382 14318 17434
rect 14330 17382 14382 17434
rect 14394 17382 14446 17434
rect 14458 17382 14510 17434
rect 14522 17382 14574 17434
rect 18705 17382 18757 17434
rect 18769 17382 18821 17434
rect 18833 17382 18885 17434
rect 18897 17382 18949 17434
rect 18961 17382 19013 17434
rect 2228 17144 2280 17196
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 3792 17144 3844 17196
rect 3976 17144 4028 17196
rect 1952 17076 2004 17128
rect 2412 17076 2464 17128
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 2044 17008 2096 17060
rect 1676 16940 1728 16992
rect 7104 16940 7156 16992
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 1860 16736 1912 16788
rect 7472 16736 7524 16788
rect 2412 16668 2464 16720
rect 2780 16668 2832 16720
rect 2964 16711 3016 16720
rect 2964 16677 2973 16711
rect 2973 16677 3007 16711
rect 3007 16677 3016 16711
rect 2964 16668 3016 16677
rect 3240 16668 3292 16720
rect 3792 16668 3844 16720
rect 940 16600 992 16652
rect 2596 16600 2648 16652
rect 3148 16600 3200 16652
rect 3976 16600 4028 16652
rect 5816 16532 5868 16584
rect 4068 16464 4120 16516
rect 4988 16464 5040 16516
rect 2780 16396 2832 16448
rect 3148 16396 3200 16448
rect 3608 16396 3660 16448
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 5644 16294 5696 16346
rect 9827 16294 9879 16346
rect 9891 16294 9943 16346
rect 9955 16294 10007 16346
rect 10019 16294 10071 16346
rect 10083 16294 10135 16346
rect 14266 16294 14318 16346
rect 14330 16294 14382 16346
rect 14394 16294 14446 16346
rect 14458 16294 14510 16346
rect 14522 16294 14574 16346
rect 18705 16294 18757 16346
rect 18769 16294 18821 16346
rect 18833 16294 18885 16346
rect 18897 16294 18949 16346
rect 18961 16294 19013 16346
rect 1584 16192 1636 16244
rect 2412 16192 2464 16244
rect 2688 16192 2740 16244
rect 5264 16192 5316 16244
rect 6184 16192 6236 16244
rect 1768 16056 1820 16108
rect 756 15920 808 15972
rect 2136 16056 2188 16108
rect 3148 16056 3200 16108
rect 2596 15988 2648 16040
rect 6276 16056 6328 16108
rect 3792 16031 3844 16040
rect 3792 15997 3801 16031
rect 3801 15997 3835 16031
rect 3835 15997 3844 16031
rect 3792 15988 3844 15997
rect 6184 15988 6236 16040
rect 2688 15920 2740 15972
rect 2872 15920 2924 15972
rect 1952 15852 2004 15904
rect 2136 15852 2188 15904
rect 2596 15852 2648 15904
rect 6460 15920 6512 15972
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 2136 15648 2188 15700
rect 2688 15648 2740 15700
rect 7472 15648 7524 15700
rect 2596 15623 2648 15632
rect 2596 15589 2605 15623
rect 2605 15589 2639 15623
rect 2639 15589 2648 15623
rect 2596 15580 2648 15589
rect 1400 15444 1452 15496
rect 4712 15444 4764 15496
rect 1952 15419 2004 15428
rect 1952 15385 1961 15419
rect 1961 15385 1995 15419
rect 1995 15385 2004 15419
rect 1952 15376 2004 15385
rect 1768 15308 1820 15360
rect 2872 15376 2924 15428
rect 5908 15444 5960 15496
rect 6184 15444 6236 15496
rect 5080 15308 5132 15360
rect 8852 15308 8904 15360
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 5644 15206 5696 15258
rect 9827 15206 9879 15258
rect 9891 15206 9943 15258
rect 9955 15206 10007 15258
rect 10019 15206 10071 15258
rect 10083 15206 10135 15258
rect 14266 15206 14318 15258
rect 14330 15206 14382 15258
rect 14394 15206 14446 15258
rect 14458 15206 14510 15258
rect 14522 15206 14574 15258
rect 18705 15206 18757 15258
rect 18769 15206 18821 15258
rect 18833 15206 18885 15258
rect 18897 15206 18949 15258
rect 18961 15206 19013 15258
rect 2320 15147 2372 15156
rect 2320 15113 2329 15147
rect 2329 15113 2363 15147
rect 2363 15113 2372 15147
rect 2320 15104 2372 15113
rect 2412 15104 2464 15156
rect 2872 15104 2924 15156
rect 5724 15104 5776 15156
rect 5908 15104 5960 15156
rect 8116 15104 8168 15156
rect 6828 15079 6880 15088
rect 6828 15045 6862 15079
rect 6862 15045 6880 15079
rect 6828 15036 6880 15045
rect 2688 14968 2740 15020
rect 6276 14968 6328 15020
rect 7932 14968 7984 15020
rect 8116 14968 8168 15020
rect 3792 14900 3844 14952
rect 3976 14900 4028 14952
rect 5816 14943 5868 14952
rect 5816 14909 5825 14943
rect 5825 14909 5859 14943
rect 5859 14909 5868 14943
rect 5816 14900 5868 14909
rect 6184 14900 6236 14952
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 4068 14560 4120 14612
rect 4252 14560 4304 14612
rect 5724 14560 5776 14612
rect 2136 14356 2188 14408
rect 3424 14356 3476 14408
rect 3976 14356 4028 14408
rect 5816 14356 5868 14408
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 6460 14399 6512 14408
rect 6460 14365 6494 14399
rect 6494 14365 6512 14399
rect 6460 14356 6512 14365
rect 1952 14288 2004 14340
rect 5264 14331 5316 14340
rect 5264 14297 5282 14331
rect 5282 14297 5316 14331
rect 5264 14288 5316 14297
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 5644 14118 5696 14170
rect 9827 14118 9879 14170
rect 9891 14118 9943 14170
rect 9955 14118 10007 14170
rect 10019 14118 10071 14170
rect 10083 14118 10135 14170
rect 14266 14118 14318 14170
rect 14330 14118 14382 14170
rect 14394 14118 14446 14170
rect 14458 14118 14510 14170
rect 14522 14118 14574 14170
rect 18705 14118 18757 14170
rect 18769 14118 18821 14170
rect 18833 14118 18885 14170
rect 18897 14118 18949 14170
rect 18961 14118 19013 14170
rect 2688 14059 2740 14068
rect 2688 14025 2690 14059
rect 2690 14025 2724 14059
rect 2724 14025 2740 14059
rect 2688 14016 2740 14025
rect 4712 14016 4764 14068
rect 5264 14016 5316 14068
rect 5908 14016 5960 14068
rect 1860 13880 1912 13932
rect 2504 13923 2556 13932
rect 2504 13889 2513 13923
rect 2513 13889 2547 13923
rect 2547 13889 2556 13923
rect 2504 13880 2556 13889
rect 2872 13880 2924 13932
rect 3056 13880 3108 13932
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 1216 13812 1268 13864
rect 4436 13880 4488 13932
rect 8760 13880 8812 13932
rect 3976 13812 4028 13864
rect 6184 13812 6236 13864
rect 6460 13812 6512 13864
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 4896 13472 4948 13524
rect 3056 13404 3108 13456
rect 4068 13404 4120 13456
rect 1952 13336 2004 13388
rect 2412 13336 2464 13388
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 2780 13268 2832 13277
rect 2872 13200 2924 13252
rect 5264 13243 5316 13252
rect 5264 13209 5273 13243
rect 5273 13209 5307 13243
rect 5307 13209 5316 13243
rect 5264 13200 5316 13209
rect 6460 13132 6512 13184
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 5644 13030 5696 13082
rect 9827 13030 9879 13082
rect 9891 13030 9943 13082
rect 9955 13030 10007 13082
rect 10019 13030 10071 13082
rect 10083 13030 10135 13082
rect 14266 13030 14318 13082
rect 14330 13030 14382 13082
rect 14394 13030 14446 13082
rect 14458 13030 14510 13082
rect 14522 13030 14574 13082
rect 18705 13030 18757 13082
rect 18769 13030 18821 13082
rect 18833 13030 18885 13082
rect 18897 13030 18949 13082
rect 18961 13030 19013 13082
rect 2136 12928 2188 12980
rect 7104 12928 7156 12980
rect 8668 12860 8720 12912
rect 2780 12792 2832 12844
rect 4068 12792 4120 12844
rect 5264 12792 5316 12844
rect 6460 12724 6512 12776
rect 2044 12699 2096 12708
rect 2044 12665 2053 12699
rect 2053 12665 2087 12699
rect 2087 12665 2096 12699
rect 2044 12656 2096 12665
rect 3608 12656 3660 12708
rect 1124 12588 1176 12640
rect 3976 12588 4028 12640
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 2872 12384 2924 12436
rect 3700 12384 3752 12436
rect 940 12316 992 12368
rect 4436 12248 4488 12300
rect 6000 12248 6052 12300
rect 6460 12248 6512 12300
rect 1952 12180 2004 12232
rect 2320 12180 2372 12232
rect 1676 12112 1728 12164
rect 2136 12112 2188 12164
rect 1032 12044 1084 12096
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 2872 12180 2924 12232
rect 2872 12044 2924 12096
rect 3516 12044 3568 12096
rect 6736 12044 6788 12096
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 5644 11942 5696 11994
rect 9827 11942 9879 11994
rect 9891 11942 9943 11994
rect 9955 11942 10007 11994
rect 10019 11942 10071 11994
rect 10083 11942 10135 11994
rect 14266 11942 14318 11994
rect 14330 11942 14382 11994
rect 14394 11942 14446 11994
rect 14458 11942 14510 11994
rect 14522 11942 14574 11994
rect 18705 11942 18757 11994
rect 18769 11942 18821 11994
rect 18833 11942 18885 11994
rect 18897 11942 18949 11994
rect 18961 11942 19013 11994
rect 2320 11840 2372 11892
rect 4712 11840 4764 11892
rect 1768 11815 1820 11824
rect 1768 11781 1777 11815
rect 1777 11781 1811 11815
rect 1811 11781 1820 11815
rect 1768 11772 1820 11781
rect 1860 11772 1912 11824
rect 2136 11815 2188 11824
rect 2136 11781 2145 11815
rect 2145 11781 2179 11815
rect 2179 11781 2188 11815
rect 2136 11772 2188 11781
rect 3976 11772 4028 11824
rect 1308 11704 1360 11756
rect 2780 11704 2832 11756
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 3516 11704 3568 11756
rect 4344 11704 4396 11756
rect 5724 11704 5776 11756
rect 6460 11704 6512 11756
rect 2412 11636 2464 11688
rect 3608 11568 3660 11620
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 1400 11296 1452 11348
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 4068 11296 4120 11348
rect 1676 11160 1728 11212
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 1952 11092 2004 11144
rect 1584 11067 1636 11076
rect 1584 11033 1593 11067
rect 1593 11033 1627 11067
rect 1627 11033 1636 11067
rect 1584 11024 1636 11033
rect 3608 11024 3660 11076
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 5644 10854 5696 10906
rect 9827 10854 9879 10906
rect 9891 10854 9943 10906
rect 9955 10854 10007 10906
rect 10019 10854 10071 10906
rect 10083 10854 10135 10906
rect 14266 10854 14318 10906
rect 14330 10854 14382 10906
rect 14394 10854 14446 10906
rect 14458 10854 14510 10906
rect 14522 10854 14574 10906
rect 18705 10854 18757 10906
rect 18769 10854 18821 10906
rect 18833 10854 18885 10906
rect 18897 10854 18949 10906
rect 18961 10854 19013 10906
rect 6368 10752 6420 10804
rect 6000 10616 6052 10668
rect 9036 10616 9088 10668
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 4620 10208 4672 10260
rect 5264 10140 5316 10192
rect 3976 10115 4028 10124
rect 3976 10081 3985 10115
rect 3985 10081 4019 10115
rect 4019 10081 4028 10115
rect 3976 10072 4028 10081
rect 940 10004 992 10056
rect 4252 10047 4304 10056
rect 4252 10013 4286 10047
rect 4286 10013 4304 10047
rect 4252 10004 4304 10013
rect 5816 9979 5868 9988
rect 5816 9945 5825 9979
rect 5825 9945 5859 9979
rect 5859 9945 5868 9979
rect 5816 9936 5868 9945
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 5644 9766 5696 9818
rect 9827 9766 9879 9818
rect 9891 9766 9943 9818
rect 9955 9766 10007 9818
rect 10019 9766 10071 9818
rect 10083 9766 10135 9818
rect 14266 9766 14318 9818
rect 14330 9766 14382 9818
rect 14394 9766 14446 9818
rect 14458 9766 14510 9818
rect 14522 9766 14574 9818
rect 18705 9766 18757 9818
rect 18769 9766 18821 9818
rect 18833 9766 18885 9818
rect 18897 9766 18949 9818
rect 18961 9766 19013 9818
rect 1768 9596 1820 9648
rect 1952 9596 2004 9648
rect 6644 9596 6696 9648
rect 8024 9460 8076 9512
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 2136 9324 2188 9376
rect 4160 9324 4212 9376
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 3148 9120 3200 9172
rect 3976 9120 4028 9172
rect 1492 9052 1544 9104
rect 2044 8984 2096 9036
rect 2504 8984 2556 9036
rect 3976 8984 4028 9036
rect 1860 8916 1912 8968
rect 1400 8848 1452 8900
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 2596 8780 2648 8832
rect 3792 8780 3844 8832
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 5644 8678 5696 8730
rect 9827 8678 9879 8730
rect 9891 8678 9943 8730
rect 9955 8678 10007 8730
rect 10019 8678 10071 8730
rect 10083 8678 10135 8730
rect 14266 8678 14318 8730
rect 14330 8678 14382 8730
rect 14394 8678 14446 8730
rect 14458 8678 14510 8730
rect 14522 8678 14574 8730
rect 18705 8678 18757 8730
rect 18769 8678 18821 8730
rect 18833 8678 18885 8730
rect 18897 8678 18949 8730
rect 18961 8678 19013 8730
rect 2780 8576 2832 8628
rect 3056 8576 3108 8628
rect 4804 8576 4856 8628
rect 2688 8551 2740 8560
rect 2688 8517 2697 8551
rect 2697 8517 2731 8551
rect 2731 8517 2740 8551
rect 2688 8508 2740 8517
rect 6552 8508 6604 8560
rect 2964 8440 3016 8492
rect 3700 8440 3752 8492
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 3792 8415 3844 8424
rect 3792 8381 3801 8415
rect 3801 8381 3835 8415
rect 3835 8381 3844 8415
rect 3792 8372 3844 8381
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 2872 7896 2924 7948
rect 756 7828 808 7880
rect 3700 7828 3752 7880
rect 1860 7692 1912 7744
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 5644 7590 5696 7642
rect 9827 7590 9879 7642
rect 9891 7590 9943 7642
rect 9955 7590 10007 7642
rect 10019 7590 10071 7642
rect 10083 7590 10135 7642
rect 14266 7590 14318 7642
rect 14330 7590 14382 7642
rect 14394 7590 14446 7642
rect 14458 7590 14510 7642
rect 14522 7590 14574 7642
rect 18705 7590 18757 7642
rect 18769 7590 18821 7642
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 7196 7488 7248 7540
rect 1308 7420 1360 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2412 7395 2464 7404
rect 2412 7361 2421 7395
rect 2421 7361 2455 7395
rect 2455 7361 2464 7395
rect 2412 7352 2464 7361
rect 8392 7420 8444 7472
rect 8208 7352 8260 7404
rect 2320 7327 2372 7336
rect 2320 7293 2329 7327
rect 2329 7293 2363 7327
rect 2363 7293 2372 7327
rect 2320 7284 2372 7293
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 6276 6944 6328 6996
rect 1860 6876 1912 6928
rect 1400 6808 1452 6860
rect 1584 6740 1636 6792
rect 2504 6808 2556 6860
rect 3792 6808 3844 6860
rect 1676 6604 1728 6656
rect 2228 6740 2280 6792
rect 2964 6740 3016 6792
rect 3884 6740 3936 6792
rect 5172 6740 5224 6792
rect 7104 6672 7156 6724
rect 8208 6672 8260 6724
rect 2688 6647 2740 6656
rect 2688 6613 2697 6647
rect 2697 6613 2731 6647
rect 2731 6613 2740 6647
rect 2688 6604 2740 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 3976 6604 4028 6656
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 5644 6502 5696 6554
rect 9827 6502 9879 6554
rect 9891 6502 9943 6554
rect 9955 6502 10007 6554
rect 10019 6502 10071 6554
rect 10083 6502 10135 6554
rect 14266 6502 14318 6554
rect 14330 6502 14382 6554
rect 14394 6502 14446 6554
rect 14458 6502 14510 6554
rect 14522 6502 14574 6554
rect 18705 6502 18757 6554
rect 18769 6502 18821 6554
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 1676 6400 1728 6452
rect 2504 6400 2556 6452
rect 4620 6443 4672 6452
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 1860 6264 1912 6316
rect 3056 6332 3108 6384
rect 7104 6332 7156 6384
rect 1952 6196 2004 6248
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6828 6307 6880 6316
rect 6828 6273 6862 6307
rect 6862 6273 6880 6307
rect 6828 6264 6880 6273
rect 7288 6400 7340 6452
rect 9680 6264 9732 6316
rect 4896 6060 4948 6112
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 2412 5856 2464 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 6828 5856 6880 5908
rect 8484 5856 8536 5908
rect 2964 5652 3016 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 940 5584 992 5636
rect 1768 5627 1820 5636
rect 1768 5593 1777 5627
rect 1777 5593 1811 5627
rect 1811 5593 1820 5627
rect 1768 5584 1820 5593
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 5644 5414 5696 5466
rect 9827 5414 9879 5466
rect 9891 5414 9943 5466
rect 9955 5414 10007 5466
rect 10019 5414 10071 5466
rect 10083 5414 10135 5466
rect 14266 5414 14318 5466
rect 14330 5414 14382 5466
rect 14394 5414 14446 5466
rect 14458 5414 14510 5466
rect 14522 5414 14574 5466
rect 18705 5414 18757 5466
rect 18769 5414 18821 5466
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 2044 5312 2096 5364
rect 3792 5312 3844 5364
rect 8116 5312 8168 5364
rect 5264 5244 5316 5296
rect 8576 5244 8628 5296
rect 1400 5176 1452 5228
rect 1860 5176 1912 5228
rect 2044 5176 2096 5228
rect 3608 5176 3660 5228
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 4988 5040 5040 5092
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 1768 4768 1820 4820
rect 3792 4632 3844 4684
rect 6552 4768 6604 4820
rect 4068 4564 4120 4616
rect 4804 4564 4856 4616
rect 6460 4607 6512 4616
rect 6460 4573 6494 4607
rect 6494 4573 6512 4607
rect 6460 4564 6512 4573
rect 7380 4496 7432 4548
rect 6000 4428 6052 4480
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 5644 4326 5696 4378
rect 9827 4326 9879 4378
rect 9891 4326 9943 4378
rect 9955 4326 10007 4378
rect 10019 4326 10071 4378
rect 10083 4326 10135 4378
rect 14266 4326 14318 4378
rect 14330 4326 14382 4378
rect 14394 4326 14446 4378
rect 14458 4326 14510 4378
rect 14522 4326 14574 4378
rect 18705 4326 18757 4378
rect 18769 4326 18821 4378
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 1124 4156 1176 4208
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2780 4156 2832 4208
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 4896 4088 4948 4140
rect 6276 4088 6328 4140
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 3056 4020 3108 4072
rect 6092 4020 6144 4072
rect 2044 3952 2096 4004
rect 2964 3952 3016 4004
rect 2596 3884 2648 3936
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 1952 3680 2004 3732
rect 6736 3680 6788 3732
rect 9128 3680 9180 3732
rect 2320 3612 2372 3664
rect 1676 3544 1728 3596
rect 3516 3544 3568 3596
rect 3792 3544 3844 3596
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 7012 3544 7064 3596
rect 4252 3519 4304 3528
rect 4252 3485 4286 3519
rect 4286 3485 4304 3519
rect 4252 3476 4304 3485
rect 4988 3476 5040 3528
rect 5816 3476 5868 3528
rect 2596 3451 2648 3460
rect 2596 3417 2605 3451
rect 2605 3417 2639 3451
rect 2639 3417 2648 3451
rect 2596 3408 2648 3417
rect 848 3340 900 3392
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 5644 3238 5696 3290
rect 9827 3238 9879 3290
rect 9891 3238 9943 3290
rect 9955 3238 10007 3290
rect 10019 3238 10071 3290
rect 10083 3238 10135 3290
rect 14266 3238 14318 3290
rect 14330 3238 14382 3290
rect 14394 3238 14446 3290
rect 14458 3238 14510 3290
rect 14522 3238 14574 3290
rect 18705 3238 18757 3290
rect 18769 3238 18821 3290
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 4160 3136 4212 3188
rect 1584 3000 1636 3052
rect 2228 3000 2280 3052
rect 3792 3000 3844 3052
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 1860 2975 1912 2984
rect 1860 2941 1869 2975
rect 1869 2941 1903 2975
rect 1903 2941 1912 2975
rect 1860 2932 1912 2941
rect 2688 2796 2740 2848
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 1216 2592 1268 2644
rect 3700 2592 3752 2644
rect 940 2456 992 2508
rect 3792 2456 3844 2508
rect 8944 2456 8996 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 5080 2388 5132 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 1952 2320 2004 2372
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 5644 2150 5696 2202
rect 9827 2150 9879 2202
rect 9891 2150 9943 2202
rect 9955 2150 10007 2202
rect 10019 2150 10071 2202
rect 10083 2150 10135 2202
rect 14266 2150 14318 2202
rect 14330 2150 14382 2202
rect 14394 2150 14446 2202
rect 14458 2150 14510 2202
rect 14522 2150 14574 2202
rect 18705 2150 18757 2202
rect 18769 2150 18821 2202
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
<< metal2 >>
rect 938 47968 994 47977
rect 938 47903 994 47912
rect 952 47190 980 47903
rect 3169 47356 3477 47365
rect 3169 47354 3175 47356
rect 3231 47354 3255 47356
rect 3311 47354 3335 47356
rect 3391 47354 3415 47356
rect 3471 47354 3477 47356
rect 3231 47302 3233 47354
rect 3413 47302 3415 47354
rect 3169 47300 3175 47302
rect 3231 47300 3255 47302
rect 3311 47300 3335 47302
rect 3391 47300 3415 47302
rect 3471 47300 3477 47302
rect 3169 47291 3477 47300
rect 7608 47356 7916 47365
rect 7608 47354 7614 47356
rect 7670 47354 7694 47356
rect 7750 47354 7774 47356
rect 7830 47354 7854 47356
rect 7910 47354 7916 47356
rect 7670 47302 7672 47354
rect 7852 47302 7854 47354
rect 7608 47300 7614 47302
rect 7670 47300 7694 47302
rect 7750 47300 7774 47302
rect 7830 47300 7854 47302
rect 7910 47300 7916 47302
rect 7608 47291 7916 47300
rect 12047 47356 12355 47365
rect 12047 47354 12053 47356
rect 12109 47354 12133 47356
rect 12189 47354 12213 47356
rect 12269 47354 12293 47356
rect 12349 47354 12355 47356
rect 12109 47302 12111 47354
rect 12291 47302 12293 47354
rect 12047 47300 12053 47302
rect 12109 47300 12133 47302
rect 12189 47300 12213 47302
rect 12269 47300 12293 47302
rect 12349 47300 12355 47302
rect 12047 47291 12355 47300
rect 16486 47356 16794 47365
rect 16486 47354 16492 47356
rect 16548 47354 16572 47356
rect 16628 47354 16652 47356
rect 16708 47354 16732 47356
rect 16788 47354 16794 47356
rect 16548 47302 16550 47354
rect 16730 47302 16732 47354
rect 16486 47300 16492 47302
rect 16548 47300 16572 47302
rect 16628 47300 16652 47302
rect 16708 47300 16732 47302
rect 16788 47300 16794 47302
rect 16486 47291 16794 47300
rect 940 47184 992 47190
rect 940 47126 992 47132
rect 1400 46980 1452 46986
rect 1400 46922 1452 46928
rect 940 44872 992 44878
rect 940 44814 992 44820
rect 952 44441 980 44814
rect 938 44432 994 44441
rect 938 44367 994 44376
rect 940 40996 992 41002
rect 940 40938 992 40944
rect 952 40905 980 40938
rect 938 40896 994 40905
rect 938 40831 994 40840
rect 940 37664 992 37670
rect 940 37606 992 37612
rect 952 37369 980 37606
rect 938 37360 994 37369
rect 938 37295 994 37304
rect 940 33924 992 33930
rect 940 33866 992 33872
rect 952 33833 980 33866
rect 938 33824 994 33833
rect 938 33759 994 33768
rect 940 30728 992 30734
rect 940 30670 992 30676
rect 952 30297 980 30670
rect 938 30288 994 30297
rect 938 30223 994 30232
rect 940 26852 992 26858
rect 940 26794 992 26800
rect 952 26761 980 26794
rect 938 26752 994 26761
rect 938 26687 994 26696
rect 1032 24132 1084 24138
rect 1032 24074 1084 24080
rect 940 23520 992 23526
rect 940 23462 992 23468
rect 952 23225 980 23462
rect 938 23216 994 23225
rect 938 23151 994 23160
rect 940 19780 992 19786
rect 940 19722 992 19728
rect 952 19689 980 19722
rect 938 19680 994 19689
rect 938 19615 994 19624
rect 940 16652 992 16658
rect 940 16594 992 16600
rect 952 16153 980 16594
rect 938 16144 994 16153
rect 938 16079 994 16088
rect 756 15972 808 15978
rect 756 15914 808 15920
rect 768 7886 796 15914
rect 938 12608 994 12617
rect 938 12543 994 12552
rect 952 12374 980 12543
rect 940 12368 992 12374
rect 940 12310 992 12316
rect 1044 12186 1072 24074
rect 1216 19848 1268 19854
rect 1216 19790 1268 19796
rect 1228 13870 1256 19790
rect 1412 15502 1440 46922
rect 5388 46812 5696 46821
rect 5388 46810 5394 46812
rect 5450 46810 5474 46812
rect 5530 46810 5554 46812
rect 5610 46810 5634 46812
rect 5690 46810 5696 46812
rect 5450 46758 5452 46810
rect 5632 46758 5634 46810
rect 5388 46756 5394 46758
rect 5450 46756 5474 46758
rect 5530 46756 5554 46758
rect 5610 46756 5634 46758
rect 5690 46756 5696 46758
rect 5388 46747 5696 46756
rect 9827 46812 10135 46821
rect 9827 46810 9833 46812
rect 9889 46810 9913 46812
rect 9969 46810 9993 46812
rect 10049 46810 10073 46812
rect 10129 46810 10135 46812
rect 9889 46758 9891 46810
rect 10071 46758 10073 46810
rect 9827 46756 9833 46758
rect 9889 46756 9913 46758
rect 9969 46756 9993 46758
rect 10049 46756 10073 46758
rect 10129 46756 10135 46758
rect 9827 46747 10135 46756
rect 14266 46812 14574 46821
rect 14266 46810 14272 46812
rect 14328 46810 14352 46812
rect 14408 46810 14432 46812
rect 14488 46810 14512 46812
rect 14568 46810 14574 46812
rect 14328 46758 14330 46810
rect 14510 46758 14512 46810
rect 14266 46756 14272 46758
rect 14328 46756 14352 46758
rect 14408 46756 14432 46758
rect 14488 46756 14512 46758
rect 14568 46756 14574 46758
rect 14266 46747 14574 46756
rect 18705 46812 19013 46821
rect 18705 46810 18711 46812
rect 18767 46810 18791 46812
rect 18847 46810 18871 46812
rect 18927 46810 18951 46812
rect 19007 46810 19013 46812
rect 18767 46758 18769 46810
rect 18949 46758 18951 46810
rect 18705 46756 18711 46758
rect 18767 46756 18791 46758
rect 18847 46756 18871 46758
rect 18927 46756 18951 46758
rect 19007 46756 19013 46758
rect 18705 46747 19013 46756
rect 3169 46268 3477 46277
rect 3169 46266 3175 46268
rect 3231 46266 3255 46268
rect 3311 46266 3335 46268
rect 3391 46266 3415 46268
rect 3471 46266 3477 46268
rect 3231 46214 3233 46266
rect 3413 46214 3415 46266
rect 3169 46212 3175 46214
rect 3231 46212 3255 46214
rect 3311 46212 3335 46214
rect 3391 46212 3415 46214
rect 3471 46212 3477 46214
rect 3169 46203 3477 46212
rect 7608 46268 7916 46277
rect 7608 46266 7614 46268
rect 7670 46266 7694 46268
rect 7750 46266 7774 46268
rect 7830 46266 7854 46268
rect 7910 46266 7916 46268
rect 7670 46214 7672 46266
rect 7852 46214 7854 46266
rect 7608 46212 7614 46214
rect 7670 46212 7694 46214
rect 7750 46212 7774 46214
rect 7830 46212 7854 46214
rect 7910 46212 7916 46214
rect 7608 46203 7916 46212
rect 12047 46268 12355 46277
rect 12047 46266 12053 46268
rect 12109 46266 12133 46268
rect 12189 46266 12213 46268
rect 12269 46266 12293 46268
rect 12349 46266 12355 46268
rect 12109 46214 12111 46266
rect 12291 46214 12293 46266
rect 12047 46212 12053 46214
rect 12109 46212 12133 46214
rect 12189 46212 12213 46214
rect 12269 46212 12293 46214
rect 12349 46212 12355 46214
rect 12047 46203 12355 46212
rect 16486 46268 16794 46277
rect 16486 46266 16492 46268
rect 16548 46266 16572 46268
rect 16628 46266 16652 46268
rect 16708 46266 16732 46268
rect 16788 46266 16794 46268
rect 16548 46214 16550 46266
rect 16730 46214 16732 46266
rect 16486 46212 16492 46214
rect 16548 46212 16572 46214
rect 16628 46212 16652 46214
rect 16708 46212 16732 46214
rect 16788 46212 16794 46214
rect 16486 46203 16794 46212
rect 5388 45724 5696 45733
rect 5388 45722 5394 45724
rect 5450 45722 5474 45724
rect 5530 45722 5554 45724
rect 5610 45722 5634 45724
rect 5690 45722 5696 45724
rect 5450 45670 5452 45722
rect 5632 45670 5634 45722
rect 5388 45668 5394 45670
rect 5450 45668 5474 45670
rect 5530 45668 5554 45670
rect 5610 45668 5634 45670
rect 5690 45668 5696 45670
rect 5388 45659 5696 45668
rect 9827 45724 10135 45733
rect 9827 45722 9833 45724
rect 9889 45722 9913 45724
rect 9969 45722 9993 45724
rect 10049 45722 10073 45724
rect 10129 45722 10135 45724
rect 9889 45670 9891 45722
rect 10071 45670 10073 45722
rect 9827 45668 9833 45670
rect 9889 45668 9913 45670
rect 9969 45668 9993 45670
rect 10049 45668 10073 45670
rect 10129 45668 10135 45670
rect 9827 45659 10135 45668
rect 14266 45724 14574 45733
rect 14266 45722 14272 45724
rect 14328 45722 14352 45724
rect 14408 45722 14432 45724
rect 14488 45722 14512 45724
rect 14568 45722 14574 45724
rect 14328 45670 14330 45722
rect 14510 45670 14512 45722
rect 14266 45668 14272 45670
rect 14328 45668 14352 45670
rect 14408 45668 14432 45670
rect 14488 45668 14512 45670
rect 14568 45668 14574 45670
rect 14266 45659 14574 45668
rect 18705 45724 19013 45733
rect 18705 45722 18711 45724
rect 18767 45722 18791 45724
rect 18847 45722 18871 45724
rect 18927 45722 18951 45724
rect 19007 45722 19013 45724
rect 18767 45670 18769 45722
rect 18949 45670 18951 45722
rect 18705 45668 18711 45670
rect 18767 45668 18791 45670
rect 18847 45668 18871 45670
rect 18927 45668 18951 45670
rect 19007 45668 19013 45670
rect 18705 45659 19013 45668
rect 3169 45180 3477 45189
rect 3169 45178 3175 45180
rect 3231 45178 3255 45180
rect 3311 45178 3335 45180
rect 3391 45178 3415 45180
rect 3471 45178 3477 45180
rect 3231 45126 3233 45178
rect 3413 45126 3415 45178
rect 3169 45124 3175 45126
rect 3231 45124 3255 45126
rect 3311 45124 3335 45126
rect 3391 45124 3415 45126
rect 3471 45124 3477 45126
rect 3169 45115 3477 45124
rect 7608 45180 7916 45189
rect 7608 45178 7614 45180
rect 7670 45178 7694 45180
rect 7750 45178 7774 45180
rect 7830 45178 7854 45180
rect 7910 45178 7916 45180
rect 7670 45126 7672 45178
rect 7852 45126 7854 45178
rect 7608 45124 7614 45126
rect 7670 45124 7694 45126
rect 7750 45124 7774 45126
rect 7830 45124 7854 45126
rect 7910 45124 7916 45126
rect 7608 45115 7916 45124
rect 12047 45180 12355 45189
rect 12047 45178 12053 45180
rect 12109 45178 12133 45180
rect 12189 45178 12213 45180
rect 12269 45178 12293 45180
rect 12349 45178 12355 45180
rect 12109 45126 12111 45178
rect 12291 45126 12293 45178
rect 12047 45124 12053 45126
rect 12109 45124 12133 45126
rect 12189 45124 12213 45126
rect 12269 45124 12293 45126
rect 12349 45124 12355 45126
rect 12047 45115 12355 45124
rect 16486 45180 16794 45189
rect 16486 45178 16492 45180
rect 16548 45178 16572 45180
rect 16628 45178 16652 45180
rect 16708 45178 16732 45180
rect 16788 45178 16794 45180
rect 16548 45126 16550 45178
rect 16730 45126 16732 45178
rect 16486 45124 16492 45126
rect 16548 45124 16572 45126
rect 16628 45124 16652 45126
rect 16708 45124 16732 45126
rect 16788 45124 16794 45126
rect 16486 45115 16794 45124
rect 5388 44636 5696 44645
rect 5388 44634 5394 44636
rect 5450 44634 5474 44636
rect 5530 44634 5554 44636
rect 5610 44634 5634 44636
rect 5690 44634 5696 44636
rect 5450 44582 5452 44634
rect 5632 44582 5634 44634
rect 5388 44580 5394 44582
rect 5450 44580 5474 44582
rect 5530 44580 5554 44582
rect 5610 44580 5634 44582
rect 5690 44580 5696 44582
rect 5388 44571 5696 44580
rect 9827 44636 10135 44645
rect 9827 44634 9833 44636
rect 9889 44634 9913 44636
rect 9969 44634 9993 44636
rect 10049 44634 10073 44636
rect 10129 44634 10135 44636
rect 9889 44582 9891 44634
rect 10071 44582 10073 44634
rect 9827 44580 9833 44582
rect 9889 44580 9913 44582
rect 9969 44580 9993 44582
rect 10049 44580 10073 44582
rect 10129 44580 10135 44582
rect 9827 44571 10135 44580
rect 14266 44636 14574 44645
rect 14266 44634 14272 44636
rect 14328 44634 14352 44636
rect 14408 44634 14432 44636
rect 14488 44634 14512 44636
rect 14568 44634 14574 44636
rect 14328 44582 14330 44634
rect 14510 44582 14512 44634
rect 14266 44580 14272 44582
rect 14328 44580 14352 44582
rect 14408 44580 14432 44582
rect 14488 44580 14512 44582
rect 14568 44580 14574 44582
rect 14266 44571 14574 44580
rect 18705 44636 19013 44645
rect 18705 44634 18711 44636
rect 18767 44634 18791 44636
rect 18847 44634 18871 44636
rect 18927 44634 18951 44636
rect 19007 44634 19013 44636
rect 18767 44582 18769 44634
rect 18949 44582 18951 44634
rect 18705 44580 18711 44582
rect 18767 44580 18791 44582
rect 18847 44580 18871 44582
rect 18927 44580 18951 44582
rect 19007 44580 19013 44582
rect 18705 44571 19013 44580
rect 3169 44092 3477 44101
rect 3169 44090 3175 44092
rect 3231 44090 3255 44092
rect 3311 44090 3335 44092
rect 3391 44090 3415 44092
rect 3471 44090 3477 44092
rect 3231 44038 3233 44090
rect 3413 44038 3415 44090
rect 3169 44036 3175 44038
rect 3231 44036 3255 44038
rect 3311 44036 3335 44038
rect 3391 44036 3415 44038
rect 3471 44036 3477 44038
rect 3169 44027 3477 44036
rect 7608 44092 7916 44101
rect 7608 44090 7614 44092
rect 7670 44090 7694 44092
rect 7750 44090 7774 44092
rect 7830 44090 7854 44092
rect 7910 44090 7916 44092
rect 7670 44038 7672 44090
rect 7852 44038 7854 44090
rect 7608 44036 7614 44038
rect 7670 44036 7694 44038
rect 7750 44036 7774 44038
rect 7830 44036 7854 44038
rect 7910 44036 7916 44038
rect 7608 44027 7916 44036
rect 12047 44092 12355 44101
rect 12047 44090 12053 44092
rect 12109 44090 12133 44092
rect 12189 44090 12213 44092
rect 12269 44090 12293 44092
rect 12349 44090 12355 44092
rect 12109 44038 12111 44090
rect 12291 44038 12293 44090
rect 12047 44036 12053 44038
rect 12109 44036 12133 44038
rect 12189 44036 12213 44038
rect 12269 44036 12293 44038
rect 12349 44036 12355 44038
rect 12047 44027 12355 44036
rect 16486 44092 16794 44101
rect 16486 44090 16492 44092
rect 16548 44090 16572 44092
rect 16628 44090 16652 44092
rect 16708 44090 16732 44092
rect 16788 44090 16794 44092
rect 16548 44038 16550 44090
rect 16730 44038 16732 44090
rect 16486 44036 16492 44038
rect 16548 44036 16572 44038
rect 16628 44036 16652 44038
rect 16708 44036 16732 44038
rect 16788 44036 16794 44038
rect 16486 44027 16794 44036
rect 5388 43548 5696 43557
rect 5388 43546 5394 43548
rect 5450 43546 5474 43548
rect 5530 43546 5554 43548
rect 5610 43546 5634 43548
rect 5690 43546 5696 43548
rect 5450 43494 5452 43546
rect 5632 43494 5634 43546
rect 5388 43492 5394 43494
rect 5450 43492 5474 43494
rect 5530 43492 5554 43494
rect 5610 43492 5634 43494
rect 5690 43492 5696 43494
rect 5388 43483 5696 43492
rect 9827 43548 10135 43557
rect 9827 43546 9833 43548
rect 9889 43546 9913 43548
rect 9969 43546 9993 43548
rect 10049 43546 10073 43548
rect 10129 43546 10135 43548
rect 9889 43494 9891 43546
rect 10071 43494 10073 43546
rect 9827 43492 9833 43494
rect 9889 43492 9913 43494
rect 9969 43492 9993 43494
rect 10049 43492 10073 43494
rect 10129 43492 10135 43494
rect 9827 43483 10135 43492
rect 14266 43548 14574 43557
rect 14266 43546 14272 43548
rect 14328 43546 14352 43548
rect 14408 43546 14432 43548
rect 14488 43546 14512 43548
rect 14568 43546 14574 43548
rect 14328 43494 14330 43546
rect 14510 43494 14512 43546
rect 14266 43492 14272 43494
rect 14328 43492 14352 43494
rect 14408 43492 14432 43494
rect 14488 43492 14512 43494
rect 14568 43492 14574 43494
rect 14266 43483 14574 43492
rect 18705 43548 19013 43557
rect 18705 43546 18711 43548
rect 18767 43546 18791 43548
rect 18847 43546 18871 43548
rect 18927 43546 18951 43548
rect 19007 43546 19013 43548
rect 18767 43494 18769 43546
rect 18949 43494 18951 43546
rect 18705 43492 18711 43494
rect 18767 43492 18791 43494
rect 18847 43492 18871 43494
rect 18927 43492 18951 43494
rect 19007 43492 19013 43494
rect 18705 43483 19013 43492
rect 3169 43004 3477 43013
rect 3169 43002 3175 43004
rect 3231 43002 3255 43004
rect 3311 43002 3335 43004
rect 3391 43002 3415 43004
rect 3471 43002 3477 43004
rect 3231 42950 3233 43002
rect 3413 42950 3415 43002
rect 3169 42948 3175 42950
rect 3231 42948 3255 42950
rect 3311 42948 3335 42950
rect 3391 42948 3415 42950
rect 3471 42948 3477 42950
rect 3169 42939 3477 42948
rect 7608 43004 7916 43013
rect 7608 43002 7614 43004
rect 7670 43002 7694 43004
rect 7750 43002 7774 43004
rect 7830 43002 7854 43004
rect 7910 43002 7916 43004
rect 7670 42950 7672 43002
rect 7852 42950 7854 43002
rect 7608 42948 7614 42950
rect 7670 42948 7694 42950
rect 7750 42948 7774 42950
rect 7830 42948 7854 42950
rect 7910 42948 7916 42950
rect 7608 42939 7916 42948
rect 12047 43004 12355 43013
rect 12047 43002 12053 43004
rect 12109 43002 12133 43004
rect 12189 43002 12213 43004
rect 12269 43002 12293 43004
rect 12349 43002 12355 43004
rect 12109 42950 12111 43002
rect 12291 42950 12293 43002
rect 12047 42948 12053 42950
rect 12109 42948 12133 42950
rect 12189 42948 12213 42950
rect 12269 42948 12293 42950
rect 12349 42948 12355 42950
rect 12047 42939 12355 42948
rect 16486 43004 16794 43013
rect 16486 43002 16492 43004
rect 16548 43002 16572 43004
rect 16628 43002 16652 43004
rect 16708 43002 16732 43004
rect 16788 43002 16794 43004
rect 16548 42950 16550 43002
rect 16730 42950 16732 43002
rect 16486 42948 16492 42950
rect 16548 42948 16572 42950
rect 16628 42948 16652 42950
rect 16708 42948 16732 42950
rect 16788 42948 16794 42950
rect 16486 42939 16794 42948
rect 5388 42460 5696 42469
rect 5388 42458 5394 42460
rect 5450 42458 5474 42460
rect 5530 42458 5554 42460
rect 5610 42458 5634 42460
rect 5690 42458 5696 42460
rect 5450 42406 5452 42458
rect 5632 42406 5634 42458
rect 5388 42404 5394 42406
rect 5450 42404 5474 42406
rect 5530 42404 5554 42406
rect 5610 42404 5634 42406
rect 5690 42404 5696 42406
rect 5388 42395 5696 42404
rect 9827 42460 10135 42469
rect 9827 42458 9833 42460
rect 9889 42458 9913 42460
rect 9969 42458 9993 42460
rect 10049 42458 10073 42460
rect 10129 42458 10135 42460
rect 9889 42406 9891 42458
rect 10071 42406 10073 42458
rect 9827 42404 9833 42406
rect 9889 42404 9913 42406
rect 9969 42404 9993 42406
rect 10049 42404 10073 42406
rect 10129 42404 10135 42406
rect 9827 42395 10135 42404
rect 14266 42460 14574 42469
rect 14266 42458 14272 42460
rect 14328 42458 14352 42460
rect 14408 42458 14432 42460
rect 14488 42458 14512 42460
rect 14568 42458 14574 42460
rect 14328 42406 14330 42458
rect 14510 42406 14512 42458
rect 14266 42404 14272 42406
rect 14328 42404 14352 42406
rect 14408 42404 14432 42406
rect 14488 42404 14512 42406
rect 14568 42404 14574 42406
rect 14266 42395 14574 42404
rect 18705 42460 19013 42469
rect 18705 42458 18711 42460
rect 18767 42458 18791 42460
rect 18847 42458 18871 42460
rect 18927 42458 18951 42460
rect 19007 42458 19013 42460
rect 18767 42406 18769 42458
rect 18949 42406 18951 42458
rect 18705 42404 18711 42406
rect 18767 42404 18791 42406
rect 18847 42404 18871 42406
rect 18927 42404 18951 42406
rect 19007 42404 19013 42406
rect 18705 42395 19013 42404
rect 3169 41916 3477 41925
rect 3169 41914 3175 41916
rect 3231 41914 3255 41916
rect 3311 41914 3335 41916
rect 3391 41914 3415 41916
rect 3471 41914 3477 41916
rect 3231 41862 3233 41914
rect 3413 41862 3415 41914
rect 3169 41860 3175 41862
rect 3231 41860 3255 41862
rect 3311 41860 3335 41862
rect 3391 41860 3415 41862
rect 3471 41860 3477 41862
rect 3169 41851 3477 41860
rect 7608 41916 7916 41925
rect 7608 41914 7614 41916
rect 7670 41914 7694 41916
rect 7750 41914 7774 41916
rect 7830 41914 7854 41916
rect 7910 41914 7916 41916
rect 7670 41862 7672 41914
rect 7852 41862 7854 41914
rect 7608 41860 7614 41862
rect 7670 41860 7694 41862
rect 7750 41860 7774 41862
rect 7830 41860 7854 41862
rect 7910 41860 7916 41862
rect 7608 41851 7916 41860
rect 12047 41916 12355 41925
rect 12047 41914 12053 41916
rect 12109 41914 12133 41916
rect 12189 41914 12213 41916
rect 12269 41914 12293 41916
rect 12349 41914 12355 41916
rect 12109 41862 12111 41914
rect 12291 41862 12293 41914
rect 12047 41860 12053 41862
rect 12109 41860 12133 41862
rect 12189 41860 12213 41862
rect 12269 41860 12293 41862
rect 12349 41860 12355 41862
rect 12047 41851 12355 41860
rect 16486 41916 16794 41925
rect 16486 41914 16492 41916
rect 16548 41914 16572 41916
rect 16628 41914 16652 41916
rect 16708 41914 16732 41916
rect 16788 41914 16794 41916
rect 16548 41862 16550 41914
rect 16730 41862 16732 41914
rect 16486 41860 16492 41862
rect 16548 41860 16572 41862
rect 16628 41860 16652 41862
rect 16708 41860 16732 41862
rect 16788 41860 16794 41862
rect 16486 41851 16794 41860
rect 5388 41372 5696 41381
rect 5388 41370 5394 41372
rect 5450 41370 5474 41372
rect 5530 41370 5554 41372
rect 5610 41370 5634 41372
rect 5690 41370 5696 41372
rect 5450 41318 5452 41370
rect 5632 41318 5634 41370
rect 5388 41316 5394 41318
rect 5450 41316 5474 41318
rect 5530 41316 5554 41318
rect 5610 41316 5634 41318
rect 5690 41316 5696 41318
rect 5388 41307 5696 41316
rect 9827 41372 10135 41381
rect 9827 41370 9833 41372
rect 9889 41370 9913 41372
rect 9969 41370 9993 41372
rect 10049 41370 10073 41372
rect 10129 41370 10135 41372
rect 9889 41318 9891 41370
rect 10071 41318 10073 41370
rect 9827 41316 9833 41318
rect 9889 41316 9913 41318
rect 9969 41316 9993 41318
rect 10049 41316 10073 41318
rect 10129 41316 10135 41318
rect 9827 41307 10135 41316
rect 14266 41372 14574 41381
rect 14266 41370 14272 41372
rect 14328 41370 14352 41372
rect 14408 41370 14432 41372
rect 14488 41370 14512 41372
rect 14568 41370 14574 41372
rect 14328 41318 14330 41370
rect 14510 41318 14512 41370
rect 14266 41316 14272 41318
rect 14328 41316 14352 41318
rect 14408 41316 14432 41318
rect 14488 41316 14512 41318
rect 14568 41316 14574 41318
rect 14266 41307 14574 41316
rect 18705 41372 19013 41381
rect 18705 41370 18711 41372
rect 18767 41370 18791 41372
rect 18847 41370 18871 41372
rect 18927 41370 18951 41372
rect 19007 41370 19013 41372
rect 18767 41318 18769 41370
rect 18949 41318 18951 41370
rect 18705 41316 18711 41318
rect 18767 41316 18791 41318
rect 18847 41316 18871 41318
rect 18927 41316 18951 41318
rect 19007 41316 19013 41318
rect 18705 41307 19013 41316
rect 2504 41132 2556 41138
rect 2504 41074 2556 41080
rect 1676 33924 1728 33930
rect 1676 33866 1728 33872
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1216 13864 1268 13870
rect 1216 13806 1268 13812
rect 1124 12640 1176 12646
rect 1124 12582 1176 12588
rect 860 12158 1072 12186
rect 756 7880 808 7886
rect 756 7822 808 7828
rect 860 3398 888 12158
rect 1032 12096 1084 12102
rect 1032 12038 1084 12044
rect 940 10056 992 10062
rect 940 9998 992 10004
rect 952 9081 980 9998
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 940 5636 992 5642
rect 940 5578 992 5584
rect 952 5545 980 5578
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 848 3392 900 3398
rect 848 3334 900 3340
rect 1044 2774 1072 12038
rect 1136 4214 1164 12582
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1320 7478 1348 11698
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1412 8906 1440 11290
rect 1504 9110 1532 19314
rect 1596 16250 1624 21830
rect 1688 16998 1716 33866
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1780 26625 1808 26930
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 1766 26616 1822 26625
rect 1766 26551 1822 26560
rect 2044 26240 2096 26246
rect 2044 26182 2096 26188
rect 2056 25226 2084 26182
rect 2148 25498 2176 26862
rect 2136 25492 2188 25498
rect 2136 25434 2188 25440
rect 2044 25220 2096 25226
rect 2044 25162 2096 25168
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 1768 22704 1820 22710
rect 1768 22646 1820 22652
rect 1780 19378 1808 22646
rect 1964 22642 1992 25094
rect 2056 24070 2084 25162
rect 2148 24206 2176 25434
rect 2228 25152 2280 25158
rect 2228 25094 2280 25100
rect 2240 24750 2268 25094
rect 2228 24744 2280 24750
rect 2228 24686 2280 24692
rect 2240 24274 2268 24686
rect 2228 24268 2280 24274
rect 2228 24210 2280 24216
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1860 22568 1912 22574
rect 1860 22510 1912 22516
rect 1872 21962 1900 22510
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1860 20800 1912 20806
rect 1860 20742 1912 20748
rect 1872 19446 1900 20742
rect 1964 19990 1992 22578
rect 2056 20942 2084 24006
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 1952 19984 2004 19990
rect 1952 19926 2004 19932
rect 1860 19440 1912 19446
rect 1860 19382 1912 19388
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1964 19310 1992 19926
rect 2042 19408 2098 19417
rect 2148 19378 2176 22374
rect 2240 21146 2268 24210
rect 2516 21570 2544 41074
rect 3169 40828 3477 40837
rect 3169 40826 3175 40828
rect 3231 40826 3255 40828
rect 3311 40826 3335 40828
rect 3391 40826 3415 40828
rect 3471 40826 3477 40828
rect 3231 40774 3233 40826
rect 3413 40774 3415 40826
rect 3169 40772 3175 40774
rect 3231 40772 3255 40774
rect 3311 40772 3335 40774
rect 3391 40772 3415 40774
rect 3471 40772 3477 40774
rect 3169 40763 3477 40772
rect 7608 40828 7916 40837
rect 7608 40826 7614 40828
rect 7670 40826 7694 40828
rect 7750 40826 7774 40828
rect 7830 40826 7854 40828
rect 7910 40826 7916 40828
rect 7670 40774 7672 40826
rect 7852 40774 7854 40826
rect 7608 40772 7614 40774
rect 7670 40772 7694 40774
rect 7750 40772 7774 40774
rect 7830 40772 7854 40774
rect 7910 40772 7916 40774
rect 7608 40763 7916 40772
rect 12047 40828 12355 40837
rect 12047 40826 12053 40828
rect 12109 40826 12133 40828
rect 12189 40826 12213 40828
rect 12269 40826 12293 40828
rect 12349 40826 12355 40828
rect 12109 40774 12111 40826
rect 12291 40774 12293 40826
rect 12047 40772 12053 40774
rect 12109 40772 12133 40774
rect 12189 40772 12213 40774
rect 12269 40772 12293 40774
rect 12349 40772 12355 40774
rect 12047 40763 12355 40772
rect 16486 40828 16794 40837
rect 16486 40826 16492 40828
rect 16548 40826 16572 40828
rect 16628 40826 16652 40828
rect 16708 40826 16732 40828
rect 16788 40826 16794 40828
rect 16548 40774 16550 40826
rect 16730 40774 16732 40826
rect 16486 40772 16492 40774
rect 16548 40772 16572 40774
rect 16628 40772 16652 40774
rect 16708 40772 16732 40774
rect 16788 40772 16794 40774
rect 16486 40763 16794 40772
rect 5388 40284 5696 40293
rect 5388 40282 5394 40284
rect 5450 40282 5474 40284
rect 5530 40282 5554 40284
rect 5610 40282 5634 40284
rect 5690 40282 5696 40284
rect 5450 40230 5452 40282
rect 5632 40230 5634 40282
rect 5388 40228 5394 40230
rect 5450 40228 5474 40230
rect 5530 40228 5554 40230
rect 5610 40228 5634 40230
rect 5690 40228 5696 40230
rect 5388 40219 5696 40228
rect 9827 40284 10135 40293
rect 9827 40282 9833 40284
rect 9889 40282 9913 40284
rect 9969 40282 9993 40284
rect 10049 40282 10073 40284
rect 10129 40282 10135 40284
rect 9889 40230 9891 40282
rect 10071 40230 10073 40282
rect 9827 40228 9833 40230
rect 9889 40228 9913 40230
rect 9969 40228 9993 40230
rect 10049 40228 10073 40230
rect 10129 40228 10135 40230
rect 9827 40219 10135 40228
rect 14266 40284 14574 40293
rect 14266 40282 14272 40284
rect 14328 40282 14352 40284
rect 14408 40282 14432 40284
rect 14488 40282 14512 40284
rect 14568 40282 14574 40284
rect 14328 40230 14330 40282
rect 14510 40230 14512 40282
rect 14266 40228 14272 40230
rect 14328 40228 14352 40230
rect 14408 40228 14432 40230
rect 14488 40228 14512 40230
rect 14568 40228 14574 40230
rect 14266 40219 14574 40228
rect 18705 40284 19013 40293
rect 18705 40282 18711 40284
rect 18767 40282 18791 40284
rect 18847 40282 18871 40284
rect 18927 40282 18951 40284
rect 19007 40282 19013 40284
rect 18767 40230 18769 40282
rect 18949 40230 18951 40282
rect 18705 40228 18711 40230
rect 18767 40228 18791 40230
rect 18847 40228 18871 40230
rect 18927 40228 18951 40230
rect 19007 40228 19013 40230
rect 18705 40219 19013 40228
rect 3169 39740 3477 39749
rect 3169 39738 3175 39740
rect 3231 39738 3255 39740
rect 3311 39738 3335 39740
rect 3391 39738 3415 39740
rect 3471 39738 3477 39740
rect 3231 39686 3233 39738
rect 3413 39686 3415 39738
rect 3169 39684 3175 39686
rect 3231 39684 3255 39686
rect 3311 39684 3335 39686
rect 3391 39684 3415 39686
rect 3471 39684 3477 39686
rect 3169 39675 3477 39684
rect 7608 39740 7916 39749
rect 7608 39738 7614 39740
rect 7670 39738 7694 39740
rect 7750 39738 7774 39740
rect 7830 39738 7854 39740
rect 7910 39738 7916 39740
rect 7670 39686 7672 39738
rect 7852 39686 7854 39738
rect 7608 39684 7614 39686
rect 7670 39684 7694 39686
rect 7750 39684 7774 39686
rect 7830 39684 7854 39686
rect 7910 39684 7916 39686
rect 7608 39675 7916 39684
rect 12047 39740 12355 39749
rect 12047 39738 12053 39740
rect 12109 39738 12133 39740
rect 12189 39738 12213 39740
rect 12269 39738 12293 39740
rect 12349 39738 12355 39740
rect 12109 39686 12111 39738
rect 12291 39686 12293 39738
rect 12047 39684 12053 39686
rect 12109 39684 12133 39686
rect 12189 39684 12213 39686
rect 12269 39684 12293 39686
rect 12349 39684 12355 39686
rect 12047 39675 12355 39684
rect 16486 39740 16794 39749
rect 16486 39738 16492 39740
rect 16548 39738 16572 39740
rect 16628 39738 16652 39740
rect 16708 39738 16732 39740
rect 16788 39738 16794 39740
rect 16548 39686 16550 39738
rect 16730 39686 16732 39738
rect 16486 39684 16492 39686
rect 16548 39684 16572 39686
rect 16628 39684 16652 39686
rect 16708 39684 16732 39686
rect 16788 39684 16794 39686
rect 16486 39675 16794 39684
rect 5388 39196 5696 39205
rect 5388 39194 5394 39196
rect 5450 39194 5474 39196
rect 5530 39194 5554 39196
rect 5610 39194 5634 39196
rect 5690 39194 5696 39196
rect 5450 39142 5452 39194
rect 5632 39142 5634 39194
rect 5388 39140 5394 39142
rect 5450 39140 5474 39142
rect 5530 39140 5554 39142
rect 5610 39140 5634 39142
rect 5690 39140 5696 39142
rect 5388 39131 5696 39140
rect 9827 39196 10135 39205
rect 9827 39194 9833 39196
rect 9889 39194 9913 39196
rect 9969 39194 9993 39196
rect 10049 39194 10073 39196
rect 10129 39194 10135 39196
rect 9889 39142 9891 39194
rect 10071 39142 10073 39194
rect 9827 39140 9833 39142
rect 9889 39140 9913 39142
rect 9969 39140 9993 39142
rect 10049 39140 10073 39142
rect 10129 39140 10135 39142
rect 9827 39131 10135 39140
rect 14266 39196 14574 39205
rect 14266 39194 14272 39196
rect 14328 39194 14352 39196
rect 14408 39194 14432 39196
rect 14488 39194 14512 39196
rect 14568 39194 14574 39196
rect 14328 39142 14330 39194
rect 14510 39142 14512 39194
rect 14266 39140 14272 39142
rect 14328 39140 14352 39142
rect 14408 39140 14432 39142
rect 14488 39140 14512 39142
rect 14568 39140 14574 39142
rect 14266 39131 14574 39140
rect 18705 39196 19013 39205
rect 18705 39194 18711 39196
rect 18767 39194 18791 39196
rect 18847 39194 18871 39196
rect 18927 39194 18951 39196
rect 19007 39194 19013 39196
rect 18767 39142 18769 39194
rect 18949 39142 18951 39194
rect 18705 39140 18711 39142
rect 18767 39140 18791 39142
rect 18847 39140 18871 39142
rect 18927 39140 18951 39142
rect 19007 39140 19013 39142
rect 18705 39131 19013 39140
rect 3169 38652 3477 38661
rect 3169 38650 3175 38652
rect 3231 38650 3255 38652
rect 3311 38650 3335 38652
rect 3391 38650 3415 38652
rect 3471 38650 3477 38652
rect 3231 38598 3233 38650
rect 3413 38598 3415 38650
rect 3169 38596 3175 38598
rect 3231 38596 3255 38598
rect 3311 38596 3335 38598
rect 3391 38596 3415 38598
rect 3471 38596 3477 38598
rect 3169 38587 3477 38596
rect 7608 38652 7916 38661
rect 7608 38650 7614 38652
rect 7670 38650 7694 38652
rect 7750 38650 7774 38652
rect 7830 38650 7854 38652
rect 7910 38650 7916 38652
rect 7670 38598 7672 38650
rect 7852 38598 7854 38650
rect 7608 38596 7614 38598
rect 7670 38596 7694 38598
rect 7750 38596 7774 38598
rect 7830 38596 7854 38598
rect 7910 38596 7916 38598
rect 7608 38587 7916 38596
rect 12047 38652 12355 38661
rect 12047 38650 12053 38652
rect 12109 38650 12133 38652
rect 12189 38650 12213 38652
rect 12269 38650 12293 38652
rect 12349 38650 12355 38652
rect 12109 38598 12111 38650
rect 12291 38598 12293 38650
rect 12047 38596 12053 38598
rect 12109 38596 12133 38598
rect 12189 38596 12213 38598
rect 12269 38596 12293 38598
rect 12349 38596 12355 38598
rect 12047 38587 12355 38596
rect 16486 38652 16794 38661
rect 16486 38650 16492 38652
rect 16548 38650 16572 38652
rect 16628 38650 16652 38652
rect 16708 38650 16732 38652
rect 16788 38650 16794 38652
rect 16548 38598 16550 38650
rect 16730 38598 16732 38650
rect 16486 38596 16492 38598
rect 16548 38596 16572 38598
rect 16628 38596 16652 38598
rect 16708 38596 16732 38598
rect 16788 38596 16794 38598
rect 16486 38587 16794 38596
rect 5388 38108 5696 38117
rect 5388 38106 5394 38108
rect 5450 38106 5474 38108
rect 5530 38106 5554 38108
rect 5610 38106 5634 38108
rect 5690 38106 5696 38108
rect 5450 38054 5452 38106
rect 5632 38054 5634 38106
rect 5388 38052 5394 38054
rect 5450 38052 5474 38054
rect 5530 38052 5554 38054
rect 5610 38052 5634 38054
rect 5690 38052 5696 38054
rect 5388 38043 5696 38052
rect 9827 38108 10135 38117
rect 9827 38106 9833 38108
rect 9889 38106 9913 38108
rect 9969 38106 9993 38108
rect 10049 38106 10073 38108
rect 10129 38106 10135 38108
rect 9889 38054 9891 38106
rect 10071 38054 10073 38106
rect 9827 38052 9833 38054
rect 9889 38052 9913 38054
rect 9969 38052 9993 38054
rect 10049 38052 10073 38054
rect 10129 38052 10135 38054
rect 9827 38043 10135 38052
rect 14266 38108 14574 38117
rect 14266 38106 14272 38108
rect 14328 38106 14352 38108
rect 14408 38106 14432 38108
rect 14488 38106 14512 38108
rect 14568 38106 14574 38108
rect 14328 38054 14330 38106
rect 14510 38054 14512 38106
rect 14266 38052 14272 38054
rect 14328 38052 14352 38054
rect 14408 38052 14432 38054
rect 14488 38052 14512 38054
rect 14568 38052 14574 38054
rect 14266 38043 14574 38052
rect 18705 38108 19013 38117
rect 18705 38106 18711 38108
rect 18767 38106 18791 38108
rect 18847 38106 18871 38108
rect 18927 38106 18951 38108
rect 19007 38106 19013 38108
rect 18767 38054 18769 38106
rect 18949 38054 18951 38106
rect 18705 38052 18711 38054
rect 18767 38052 18791 38054
rect 18847 38052 18871 38054
rect 18927 38052 18951 38054
rect 19007 38052 19013 38054
rect 18705 38043 19013 38052
rect 3169 37564 3477 37573
rect 3169 37562 3175 37564
rect 3231 37562 3255 37564
rect 3311 37562 3335 37564
rect 3391 37562 3415 37564
rect 3471 37562 3477 37564
rect 3231 37510 3233 37562
rect 3413 37510 3415 37562
rect 3169 37508 3175 37510
rect 3231 37508 3255 37510
rect 3311 37508 3335 37510
rect 3391 37508 3415 37510
rect 3471 37508 3477 37510
rect 3169 37499 3477 37508
rect 7608 37564 7916 37573
rect 7608 37562 7614 37564
rect 7670 37562 7694 37564
rect 7750 37562 7774 37564
rect 7830 37562 7854 37564
rect 7910 37562 7916 37564
rect 7670 37510 7672 37562
rect 7852 37510 7854 37562
rect 7608 37508 7614 37510
rect 7670 37508 7694 37510
rect 7750 37508 7774 37510
rect 7830 37508 7854 37510
rect 7910 37508 7916 37510
rect 7608 37499 7916 37508
rect 12047 37564 12355 37573
rect 12047 37562 12053 37564
rect 12109 37562 12133 37564
rect 12189 37562 12213 37564
rect 12269 37562 12293 37564
rect 12349 37562 12355 37564
rect 12109 37510 12111 37562
rect 12291 37510 12293 37562
rect 12047 37508 12053 37510
rect 12109 37508 12133 37510
rect 12189 37508 12213 37510
rect 12269 37508 12293 37510
rect 12349 37508 12355 37510
rect 12047 37499 12355 37508
rect 16486 37564 16794 37573
rect 16486 37562 16492 37564
rect 16548 37562 16572 37564
rect 16628 37562 16652 37564
rect 16708 37562 16732 37564
rect 16788 37562 16794 37564
rect 16548 37510 16550 37562
rect 16730 37510 16732 37562
rect 16486 37508 16492 37510
rect 16548 37508 16572 37510
rect 16628 37508 16652 37510
rect 16708 37508 16732 37510
rect 16788 37508 16794 37510
rect 16486 37499 16794 37508
rect 5388 37020 5696 37029
rect 5388 37018 5394 37020
rect 5450 37018 5474 37020
rect 5530 37018 5554 37020
rect 5610 37018 5634 37020
rect 5690 37018 5696 37020
rect 5450 36966 5452 37018
rect 5632 36966 5634 37018
rect 5388 36964 5394 36966
rect 5450 36964 5474 36966
rect 5530 36964 5554 36966
rect 5610 36964 5634 36966
rect 5690 36964 5696 36966
rect 5388 36955 5696 36964
rect 9827 37020 10135 37029
rect 9827 37018 9833 37020
rect 9889 37018 9913 37020
rect 9969 37018 9993 37020
rect 10049 37018 10073 37020
rect 10129 37018 10135 37020
rect 9889 36966 9891 37018
rect 10071 36966 10073 37018
rect 9827 36964 9833 36966
rect 9889 36964 9913 36966
rect 9969 36964 9993 36966
rect 10049 36964 10073 36966
rect 10129 36964 10135 36966
rect 9827 36955 10135 36964
rect 14266 37020 14574 37029
rect 14266 37018 14272 37020
rect 14328 37018 14352 37020
rect 14408 37018 14432 37020
rect 14488 37018 14512 37020
rect 14568 37018 14574 37020
rect 14328 36966 14330 37018
rect 14510 36966 14512 37018
rect 14266 36964 14272 36966
rect 14328 36964 14352 36966
rect 14408 36964 14432 36966
rect 14488 36964 14512 36966
rect 14568 36964 14574 36966
rect 14266 36955 14574 36964
rect 18705 37020 19013 37029
rect 18705 37018 18711 37020
rect 18767 37018 18791 37020
rect 18847 37018 18871 37020
rect 18927 37018 18951 37020
rect 19007 37018 19013 37020
rect 18767 36966 18769 37018
rect 18949 36966 18951 37018
rect 18705 36964 18711 36966
rect 18767 36964 18791 36966
rect 18847 36964 18871 36966
rect 18927 36964 18951 36966
rect 19007 36964 19013 36966
rect 18705 36955 19013 36964
rect 3169 36476 3477 36485
rect 3169 36474 3175 36476
rect 3231 36474 3255 36476
rect 3311 36474 3335 36476
rect 3391 36474 3415 36476
rect 3471 36474 3477 36476
rect 3231 36422 3233 36474
rect 3413 36422 3415 36474
rect 3169 36420 3175 36422
rect 3231 36420 3255 36422
rect 3311 36420 3335 36422
rect 3391 36420 3415 36422
rect 3471 36420 3477 36422
rect 3169 36411 3477 36420
rect 7608 36476 7916 36485
rect 7608 36474 7614 36476
rect 7670 36474 7694 36476
rect 7750 36474 7774 36476
rect 7830 36474 7854 36476
rect 7910 36474 7916 36476
rect 7670 36422 7672 36474
rect 7852 36422 7854 36474
rect 7608 36420 7614 36422
rect 7670 36420 7694 36422
rect 7750 36420 7774 36422
rect 7830 36420 7854 36422
rect 7910 36420 7916 36422
rect 7608 36411 7916 36420
rect 12047 36476 12355 36485
rect 12047 36474 12053 36476
rect 12109 36474 12133 36476
rect 12189 36474 12213 36476
rect 12269 36474 12293 36476
rect 12349 36474 12355 36476
rect 12109 36422 12111 36474
rect 12291 36422 12293 36474
rect 12047 36420 12053 36422
rect 12109 36420 12133 36422
rect 12189 36420 12213 36422
rect 12269 36420 12293 36422
rect 12349 36420 12355 36422
rect 12047 36411 12355 36420
rect 16486 36476 16794 36485
rect 16486 36474 16492 36476
rect 16548 36474 16572 36476
rect 16628 36474 16652 36476
rect 16708 36474 16732 36476
rect 16788 36474 16794 36476
rect 16548 36422 16550 36474
rect 16730 36422 16732 36474
rect 16486 36420 16492 36422
rect 16548 36420 16572 36422
rect 16628 36420 16652 36422
rect 16708 36420 16732 36422
rect 16788 36420 16794 36422
rect 16486 36411 16794 36420
rect 7288 36236 7340 36242
rect 7288 36178 7340 36184
rect 7196 36168 7248 36174
rect 7196 36110 7248 36116
rect 4620 36100 4672 36106
rect 4620 36042 4672 36048
rect 6920 36100 6972 36106
rect 6920 36042 6972 36048
rect 4632 35698 4660 36042
rect 5388 35932 5696 35941
rect 5388 35930 5394 35932
rect 5450 35930 5474 35932
rect 5530 35930 5554 35932
rect 5610 35930 5634 35932
rect 5690 35930 5696 35932
rect 5450 35878 5452 35930
rect 5632 35878 5634 35930
rect 5388 35876 5394 35878
rect 5450 35876 5474 35878
rect 5530 35876 5554 35878
rect 5610 35876 5634 35878
rect 5690 35876 5696 35878
rect 5388 35867 5696 35876
rect 4620 35692 4672 35698
rect 4620 35634 4672 35640
rect 6184 35692 6236 35698
rect 6184 35634 6236 35640
rect 3169 35388 3477 35397
rect 3169 35386 3175 35388
rect 3231 35386 3255 35388
rect 3311 35386 3335 35388
rect 3391 35386 3415 35388
rect 3471 35386 3477 35388
rect 3231 35334 3233 35386
rect 3413 35334 3415 35386
rect 3169 35332 3175 35334
rect 3231 35332 3255 35334
rect 3311 35332 3335 35334
rect 3391 35332 3415 35334
rect 3471 35332 3477 35334
rect 3169 35323 3477 35332
rect 3169 34300 3477 34309
rect 3169 34298 3175 34300
rect 3231 34298 3255 34300
rect 3311 34298 3335 34300
rect 3391 34298 3415 34300
rect 3471 34298 3477 34300
rect 3231 34246 3233 34298
rect 3413 34246 3415 34298
rect 3169 34244 3175 34246
rect 3231 34244 3255 34246
rect 3311 34244 3335 34246
rect 3391 34244 3415 34246
rect 3471 34244 3477 34246
rect 3169 34235 3477 34244
rect 3169 33212 3477 33221
rect 3169 33210 3175 33212
rect 3231 33210 3255 33212
rect 3311 33210 3335 33212
rect 3391 33210 3415 33212
rect 3471 33210 3477 33212
rect 3231 33158 3233 33210
rect 3413 33158 3415 33210
rect 3169 33156 3175 33158
rect 3231 33156 3255 33158
rect 3311 33156 3335 33158
rect 3391 33156 3415 33158
rect 3471 33156 3477 33158
rect 3169 33147 3477 33156
rect 4632 32434 4660 35634
rect 5264 35488 5316 35494
rect 5264 35430 5316 35436
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 5172 32428 5224 32434
rect 5172 32370 5224 32376
rect 3169 32124 3477 32133
rect 3169 32122 3175 32124
rect 3231 32122 3255 32124
rect 3311 32122 3335 32124
rect 3391 32122 3415 32124
rect 3471 32122 3477 32124
rect 3231 32070 3233 32122
rect 3413 32070 3415 32122
rect 3169 32068 3175 32070
rect 3231 32068 3255 32070
rect 3311 32068 3335 32070
rect 3391 32068 3415 32070
rect 3471 32068 3477 32070
rect 3169 32059 3477 32068
rect 4712 31748 4764 31754
rect 4712 31690 4764 31696
rect 3169 31036 3477 31045
rect 3169 31034 3175 31036
rect 3231 31034 3255 31036
rect 3311 31034 3335 31036
rect 3391 31034 3415 31036
rect 3471 31034 3477 31036
rect 3231 30982 3233 31034
rect 3413 30982 3415 31034
rect 3169 30980 3175 30982
rect 3231 30980 3255 30982
rect 3311 30980 3335 30982
rect 3391 30980 3415 30982
rect 3471 30980 3477 30982
rect 3169 30971 3477 30980
rect 4724 30433 4752 31690
rect 5184 31278 5212 32370
rect 5276 31822 5304 35430
rect 6092 35080 6144 35086
rect 6092 35022 6144 35028
rect 5388 34844 5696 34853
rect 5388 34842 5394 34844
rect 5450 34842 5474 34844
rect 5530 34842 5554 34844
rect 5610 34842 5634 34844
rect 5690 34842 5696 34844
rect 5450 34790 5452 34842
rect 5632 34790 5634 34842
rect 5388 34788 5394 34790
rect 5450 34788 5474 34790
rect 5530 34788 5554 34790
rect 5610 34788 5634 34790
rect 5690 34788 5696 34790
rect 5388 34779 5696 34788
rect 5724 34060 5776 34066
rect 5724 34002 5776 34008
rect 5388 33756 5696 33765
rect 5388 33754 5394 33756
rect 5450 33754 5474 33756
rect 5530 33754 5554 33756
rect 5610 33754 5634 33756
rect 5690 33754 5696 33756
rect 5450 33702 5452 33754
rect 5632 33702 5634 33754
rect 5388 33700 5394 33702
rect 5450 33700 5474 33702
rect 5530 33700 5554 33702
rect 5610 33700 5634 33702
rect 5690 33700 5696 33702
rect 5388 33691 5696 33700
rect 5388 32668 5696 32677
rect 5388 32666 5394 32668
rect 5450 32666 5474 32668
rect 5530 32666 5554 32668
rect 5610 32666 5634 32668
rect 5690 32666 5696 32668
rect 5450 32614 5452 32666
rect 5632 32614 5634 32666
rect 5388 32612 5394 32614
rect 5450 32612 5474 32614
rect 5530 32612 5554 32614
rect 5610 32612 5634 32614
rect 5690 32612 5696 32614
rect 5388 32603 5696 32612
rect 5736 32502 5764 34002
rect 6104 33046 6132 35022
rect 6196 34406 6224 35634
rect 6932 35086 6960 36042
rect 6920 35080 6972 35086
rect 6920 35022 6972 35028
rect 6368 34944 6420 34950
rect 6368 34886 6420 34892
rect 6184 34400 6236 34406
rect 6184 34342 6236 34348
rect 6196 34066 6224 34342
rect 6380 34202 6408 34886
rect 6932 34678 6960 35022
rect 6920 34672 6972 34678
rect 6920 34614 6972 34620
rect 6460 34604 6512 34610
rect 6460 34546 6512 34552
rect 6368 34196 6420 34202
rect 6368 34138 6420 34144
rect 6184 34060 6236 34066
rect 6184 34002 6236 34008
rect 6092 33040 6144 33046
rect 6092 32982 6144 32988
rect 6184 33040 6236 33046
rect 6184 32982 6236 32988
rect 5724 32496 5776 32502
rect 5724 32438 5776 32444
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5388 31580 5696 31589
rect 5388 31578 5394 31580
rect 5450 31578 5474 31580
rect 5530 31578 5554 31580
rect 5610 31578 5634 31580
rect 5690 31578 5696 31580
rect 5450 31526 5452 31578
rect 5632 31526 5634 31578
rect 5388 31524 5394 31526
rect 5450 31524 5474 31526
rect 5530 31524 5554 31526
rect 5610 31524 5634 31526
rect 5690 31524 5696 31526
rect 5388 31515 5696 31524
rect 5632 31340 5684 31346
rect 5632 31282 5684 31288
rect 5172 31272 5224 31278
rect 5172 31214 5224 31220
rect 5644 30682 5672 31282
rect 5736 30802 5764 32438
rect 6104 32298 6132 32982
rect 6196 32910 6224 32982
rect 6184 32904 6236 32910
rect 6184 32846 6236 32852
rect 6092 32292 6144 32298
rect 6092 32234 6144 32240
rect 5908 31816 5960 31822
rect 5908 31758 5960 31764
rect 5920 31482 5948 31758
rect 5908 31476 5960 31482
rect 5908 31418 5960 31424
rect 6000 31340 6052 31346
rect 6000 31282 6052 31288
rect 5724 30796 5776 30802
rect 5724 30738 5776 30744
rect 6012 30734 6040 31282
rect 6000 30728 6052 30734
rect 5644 30654 5764 30682
rect 6000 30670 6052 30676
rect 5388 30492 5696 30501
rect 5388 30490 5394 30492
rect 5450 30490 5474 30492
rect 5530 30490 5554 30492
rect 5610 30490 5634 30492
rect 5690 30490 5696 30492
rect 5450 30438 5452 30490
rect 5632 30438 5634 30490
rect 5388 30436 5394 30438
rect 5450 30436 5474 30438
rect 5530 30436 5554 30438
rect 5610 30436 5634 30438
rect 5690 30436 5696 30438
rect 4710 30424 4766 30433
rect 5388 30427 5696 30436
rect 4710 30359 4766 30368
rect 3169 29948 3477 29957
rect 3169 29946 3175 29948
rect 3231 29946 3255 29948
rect 3311 29946 3335 29948
rect 3391 29946 3415 29948
rect 3471 29946 3477 29948
rect 3231 29894 3233 29946
rect 3413 29894 3415 29946
rect 3169 29892 3175 29894
rect 3231 29892 3255 29894
rect 3311 29892 3335 29894
rect 3391 29892 3415 29894
rect 3471 29892 3477 29894
rect 3169 29883 3477 29892
rect 5736 29850 5764 30654
rect 6012 30598 6040 30670
rect 6000 30592 6052 30598
rect 6000 30534 6052 30540
rect 5724 29844 5776 29850
rect 5724 29786 5776 29792
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4804 29504 4856 29510
rect 4804 29446 4856 29452
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 4528 29164 4580 29170
rect 4528 29106 4580 29112
rect 3169 28860 3477 28869
rect 3169 28858 3175 28860
rect 3231 28858 3255 28860
rect 3311 28858 3335 28860
rect 3391 28858 3415 28860
rect 3471 28858 3477 28860
rect 3231 28806 3233 28858
rect 3413 28806 3415 28858
rect 3169 28804 3175 28806
rect 3231 28804 3255 28806
rect 3311 28804 3335 28806
rect 3391 28804 3415 28806
rect 3471 28804 3477 28806
rect 3169 28795 3477 28804
rect 4160 28756 4212 28762
rect 4160 28698 4212 28704
rect 4068 28552 4120 28558
rect 4068 28494 4120 28500
rect 3792 28484 3844 28490
rect 3792 28426 3844 28432
rect 3169 27772 3477 27781
rect 3169 27770 3175 27772
rect 3231 27770 3255 27772
rect 3311 27770 3335 27772
rect 3391 27770 3415 27772
rect 3471 27770 3477 27772
rect 3231 27718 3233 27770
rect 3413 27718 3415 27770
rect 3169 27716 3175 27718
rect 3231 27716 3255 27718
rect 3311 27716 3335 27718
rect 3391 27716 3415 27718
rect 3471 27716 3477 27718
rect 3169 27707 3477 27716
rect 3608 27532 3660 27538
rect 3608 27474 3660 27480
rect 3620 27130 3648 27474
rect 3804 27470 3832 28426
rect 3976 28416 4028 28422
rect 3976 28358 4028 28364
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 3608 27124 3660 27130
rect 3608 27066 3660 27072
rect 2872 27056 2924 27062
rect 2872 26998 2924 27004
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 2608 22710 2636 26386
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2596 22704 2648 22710
rect 2596 22646 2648 22652
rect 2516 21542 2636 21570
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2240 19378 2268 20878
rect 2042 19343 2044 19352
rect 2096 19343 2098 19352
rect 2136 19372 2188 19378
rect 2044 19314 2096 19320
rect 2136 19314 2188 19320
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2332 18222 2360 18702
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1872 16794 1900 17818
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1964 16574 1992 17070
rect 2044 17060 2096 17066
rect 2044 17002 2096 17008
rect 1872 16546 1992 16574
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1780 15366 1808 16050
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1872 15314 1900 16546
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1964 15434 1992 15846
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 11218 1716 12106
rect 1780 11830 1808 15302
rect 1872 15286 1992 15314
rect 1964 14346 1992 15286
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1872 11830 1900 13874
rect 1964 13394 1992 14282
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 2056 12714 2084 17002
rect 2148 16114 2176 17478
rect 2240 17202 2268 17614
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2148 15706 2176 15846
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2148 14414 2176 15642
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2148 12986 2176 14350
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1780 11354 1808 11766
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1688 11098 1716 11154
rect 1964 11150 1992 12174
rect 2148 12170 2176 12922
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2240 11880 2268 17138
rect 2332 15162 2360 18158
rect 2424 17678 2452 18226
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2424 17134 2452 17614
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 2424 16250 2452 16662
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2424 15162 2452 16186
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2424 15042 2452 15098
rect 2332 15014 2452 15042
rect 2332 12238 2360 15014
rect 2516 13938 2544 18022
rect 2608 17882 2636 21542
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2608 16658 2636 17478
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2700 16250 2728 24550
rect 2780 21956 2832 21962
rect 2780 21898 2832 21904
rect 2792 21010 2820 21898
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2792 19786 2820 20946
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2884 18850 2912 26998
rect 3169 26684 3477 26693
rect 3169 26682 3175 26684
rect 3231 26682 3255 26684
rect 3311 26682 3335 26684
rect 3391 26682 3415 26684
rect 3471 26682 3477 26684
rect 3231 26630 3233 26682
rect 3413 26630 3415 26682
rect 3169 26628 3175 26630
rect 3231 26628 3255 26630
rect 3311 26628 3335 26630
rect 3391 26628 3415 26630
rect 3471 26628 3477 26630
rect 3169 26619 3477 26628
rect 3169 25596 3477 25605
rect 3169 25594 3175 25596
rect 3231 25594 3255 25596
rect 3311 25594 3335 25596
rect 3391 25594 3415 25596
rect 3471 25594 3477 25596
rect 3231 25542 3233 25594
rect 3413 25542 3415 25594
rect 3169 25540 3175 25542
rect 3231 25540 3255 25542
rect 3311 25540 3335 25542
rect 3391 25540 3415 25542
rect 3471 25540 3477 25542
rect 3169 25531 3477 25540
rect 3620 25294 3648 27066
rect 3608 25288 3660 25294
rect 3608 25230 3660 25236
rect 3169 24508 3477 24517
rect 3169 24506 3175 24508
rect 3231 24506 3255 24508
rect 3311 24506 3335 24508
rect 3391 24506 3415 24508
rect 3471 24506 3477 24508
rect 3231 24454 3233 24506
rect 3413 24454 3415 24506
rect 3169 24452 3175 24454
rect 3231 24452 3255 24454
rect 3311 24452 3335 24454
rect 3391 24452 3415 24454
rect 3471 24452 3477 24454
rect 3169 24443 3477 24452
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 2976 20058 3004 24006
rect 3169 23420 3477 23429
rect 3169 23418 3175 23420
rect 3231 23418 3255 23420
rect 3311 23418 3335 23420
rect 3391 23418 3415 23420
rect 3471 23418 3477 23420
rect 3231 23366 3233 23418
rect 3413 23366 3415 23418
rect 3169 23364 3175 23366
rect 3231 23364 3255 23366
rect 3311 23364 3335 23366
rect 3391 23364 3415 23366
rect 3471 23364 3477 23366
rect 3169 23355 3477 23364
rect 3169 22332 3477 22341
rect 3169 22330 3175 22332
rect 3231 22330 3255 22332
rect 3311 22330 3335 22332
rect 3391 22330 3415 22332
rect 3471 22330 3477 22332
rect 3231 22278 3233 22330
rect 3413 22278 3415 22330
rect 3169 22276 3175 22278
rect 3231 22276 3255 22278
rect 3311 22276 3335 22278
rect 3391 22276 3415 22278
rect 3471 22276 3477 22278
rect 3169 22267 3477 22276
rect 3169 21244 3477 21253
rect 3169 21242 3175 21244
rect 3231 21242 3255 21244
rect 3311 21242 3335 21244
rect 3391 21242 3415 21244
rect 3471 21242 3477 21244
rect 3231 21190 3233 21242
rect 3413 21190 3415 21242
rect 3169 21188 3175 21190
rect 3231 21188 3255 21190
rect 3311 21188 3335 21190
rect 3391 21188 3415 21190
rect 3471 21188 3477 21190
rect 3169 21179 3477 21188
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 3068 20398 3096 20810
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3160 20466 3188 20742
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3068 18970 3096 20334
rect 3712 20262 3740 20878
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3169 20156 3477 20165
rect 3169 20154 3175 20156
rect 3231 20154 3255 20156
rect 3311 20154 3335 20156
rect 3391 20154 3415 20156
rect 3471 20154 3477 20156
rect 3231 20102 3233 20154
rect 3413 20102 3415 20154
rect 3169 20100 3175 20102
rect 3231 20100 3255 20102
rect 3311 20100 3335 20102
rect 3391 20100 3415 20102
rect 3471 20100 3477 20102
rect 3169 20091 3477 20100
rect 3169 19068 3477 19077
rect 3169 19066 3175 19068
rect 3231 19066 3255 19068
rect 3311 19066 3335 19068
rect 3391 19066 3415 19068
rect 3471 19066 3477 19068
rect 3231 19014 3233 19066
rect 3413 19014 3415 19066
rect 3169 19012 3175 19014
rect 3231 19012 3255 19014
rect 3311 19012 3335 19014
rect 3391 19012 3415 19014
rect 3471 19012 3477 19014
rect 3169 19003 3477 19012
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3712 18850 3740 20198
rect 3804 18970 3832 27406
rect 3988 20874 4016 28358
rect 4080 27470 4108 28494
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 4080 27062 4108 27406
rect 4172 27130 4200 28698
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4264 27713 4292 28358
rect 4250 27704 4306 27713
rect 4250 27639 4306 27648
rect 4252 27600 4304 27606
rect 4252 27542 4304 27548
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4080 24954 4108 25230
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 4080 23866 4108 24890
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 4172 24410 4200 24550
rect 4160 24404 4212 24410
rect 4160 24346 4212 24352
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4264 23730 4292 27542
rect 4436 27464 4488 27470
rect 4436 27406 4488 27412
rect 4344 26988 4396 26994
rect 4344 26930 4396 26936
rect 4356 26450 4384 26930
rect 4448 26586 4476 27406
rect 4540 26586 4568 29106
rect 4632 28694 4660 29446
rect 4816 29102 4844 29446
rect 4908 29238 4936 29446
rect 4896 29232 4948 29238
rect 4896 29174 4948 29180
rect 5000 29102 5028 29582
rect 5080 29572 5132 29578
rect 5080 29514 5132 29520
rect 5092 29102 5120 29514
rect 5388 29404 5696 29413
rect 5388 29402 5394 29404
rect 5450 29402 5474 29404
rect 5530 29402 5554 29404
rect 5610 29402 5634 29404
rect 5690 29402 5696 29404
rect 5450 29350 5452 29402
rect 5632 29350 5634 29402
rect 5388 29348 5394 29350
rect 5450 29348 5474 29350
rect 5530 29348 5554 29350
rect 5610 29348 5634 29350
rect 5690 29348 5696 29350
rect 5388 29339 5696 29348
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4988 29096 5040 29102
rect 4988 29038 5040 29044
rect 5080 29096 5132 29102
rect 5080 29038 5132 29044
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4620 28688 4672 28694
rect 4620 28630 4672 28636
rect 4724 28490 4752 28902
rect 4712 28484 4764 28490
rect 4712 28426 4764 28432
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4436 26580 4488 26586
rect 4436 26522 4488 26528
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 4448 25974 4476 26522
rect 4436 25968 4488 25974
rect 4436 25910 4488 25916
rect 4344 25900 4396 25906
rect 4344 25842 4396 25848
rect 4356 24070 4384 25842
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4080 23497 4108 23666
rect 4252 23588 4304 23594
rect 4252 23530 4304 23536
rect 4066 23488 4122 23497
rect 4066 23423 4122 23432
rect 4080 22710 4108 23423
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 3976 19780 4028 19786
rect 3976 19722 4028 19728
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 2780 18828 2832 18834
rect 2884 18822 3556 18850
rect 3712 18822 3832 18850
rect 2780 18770 2832 18776
rect 2792 16726 2820 18770
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3252 18290 3280 18702
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2884 17202 2912 18090
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2976 16810 3004 17818
rect 2884 16782 3004 16810
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2608 15910 2636 15982
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2700 15706 2728 15914
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2608 13954 2636 15574
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2700 14074 2728 14962
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2504 13932 2556 13938
rect 2608 13926 2728 13954
rect 2504 13874 2556 13880
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2320 11892 2372 11898
rect 2240 11852 2320 11880
rect 2320 11834 2372 11840
rect 2136 11824 2188 11830
rect 2188 11772 2268 11778
rect 2136 11766 2268 11772
rect 2148 11750 2268 11766
rect 1952 11144 2004 11150
rect 1584 11076 1636 11082
rect 1688 11070 1808 11098
rect 1952 11086 2004 11092
rect 1584 11018 1636 11024
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 1400 8900 1452 8906
rect 1400 8842 1452 8848
rect 1308 7472 1360 7478
rect 1308 7414 1360 7420
rect 1412 6866 1440 8842
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 5234 1440 6802
rect 1596 6798 1624 11018
rect 1780 9654 1808 11070
rect 1964 9738 1992 11086
rect 1964 9710 2084 9738
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1780 6746 1808 9590
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 7750 1900 8910
rect 1964 8838 1992 9590
rect 2056 9042 2084 9710
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 6934 1900 7686
rect 1860 6928 1912 6934
rect 1860 6870 1912 6876
rect 1780 6718 1900 6746
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 6458 1716 6598
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1688 4706 1716 6394
rect 1872 6322 1900 6718
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1872 6100 1900 6258
rect 1964 6254 1992 8774
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1872 6072 1992 6100
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1780 4826 1808 5578
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1688 4678 1808 4706
rect 1124 4208 1176 4214
rect 1124 4150 1176 4156
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3602 1716 4082
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1044 2746 1256 2774
rect 1228 2650 1256 2746
rect 1216 2644 1268 2650
rect 1216 2586 1268 2592
rect 940 2508 992 2514
rect 940 2450 992 2456
rect 952 2009 980 2450
rect 1596 2446 1624 2994
rect 1780 2990 1808 4678
rect 1872 2990 1900 5170
rect 1964 5030 1992 6072
rect 2056 5370 2084 7142
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1964 3738 1992 4966
rect 2056 4010 2084 5170
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2148 3194 2176 9318
rect 2240 7410 2268 11750
rect 2332 8430 2360 11834
rect 2424 11694 2452 13330
rect 2700 12238 2728 13926
rect 2792 13920 2820 16390
rect 2884 15978 2912 16782
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2884 15162 2912 15370
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2872 13932 2924 13938
rect 2792 13892 2872 13920
rect 2872 13874 2924 13880
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12850 2820 13262
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2778 12744 2834 12753
rect 2778 12679 2834 12688
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2792 11762 2820 12679
rect 2884 12442 2912 13194
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 12102 2912 12174
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2332 7342 2360 8366
rect 2424 7410 2452 11630
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2240 3058 2268 6734
rect 2332 3670 2360 7278
rect 2516 6866 2544 8978
rect 2596 8832 2648 8838
rect 2792 8786 2820 9687
rect 2596 8774 2648 8780
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 6458 2544 6802
rect 2608 6644 2636 8774
rect 2700 8758 2820 8786
rect 2700 8566 2728 8758
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2700 6769 2728 8502
rect 2686 6760 2742 6769
rect 2686 6695 2742 6704
rect 2688 6656 2740 6662
rect 2608 6616 2688 6644
rect 2688 6598 2740 6604
rect 2594 6488 2650 6497
rect 2504 6452 2556 6458
rect 2594 6423 2650 6432
rect 2504 6394 2556 6400
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2424 5914 2452 6258
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2608 4078 2636 6423
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2608 3466 2636 3878
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1860 2984 1912 2990
rect 1912 2932 1992 2938
rect 1860 2926 1992 2932
rect 1780 2774 1808 2926
rect 1872 2910 1992 2926
rect 1780 2746 1900 2774
rect 1872 2446 1900 2746
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1964 2378 1992 2910
rect 2700 2854 2728 6598
rect 2792 4214 2820 8570
rect 2884 7954 2912 12038
rect 2976 11762 3004 16662
rect 3068 13938 3096 18022
rect 3169 17980 3477 17989
rect 3169 17978 3175 17980
rect 3231 17978 3255 17980
rect 3311 17978 3335 17980
rect 3391 17978 3415 17980
rect 3471 17978 3477 17980
rect 3231 17926 3233 17978
rect 3413 17926 3415 17978
rect 3169 17924 3175 17926
rect 3231 17924 3255 17926
rect 3311 17924 3335 17926
rect 3391 17924 3415 17926
rect 3471 17924 3477 17926
rect 3169 17915 3477 17924
rect 3528 17882 3556 18822
rect 3608 18692 3660 18698
rect 3608 18634 3660 18640
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 3240 16720 3292 16726
rect 3146 16688 3202 16697
rect 3240 16662 3292 16668
rect 3146 16623 3148 16632
rect 3200 16623 3202 16632
rect 3148 16594 3200 16600
rect 3252 16538 3280 16662
rect 3160 16510 3280 16538
rect 3160 16454 3188 16510
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3160 16114 3188 16390
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 13938 3464 14350
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 3068 8634 3096 13398
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 3528 12102 3556 17614
rect 3620 16454 3648 18634
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3620 12889 3648 16390
rect 3712 14770 3740 17546
rect 3804 17202 3832 18822
rect 3884 17740 3936 17746
rect 3884 17682 3936 17688
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3804 16726 3832 17138
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 14958 3832 15982
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3712 14742 3832 14770
rect 3606 12880 3662 12889
rect 3606 12815 3662 12824
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3620 11914 3648 12650
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3528 11886 3648 11914
rect 3528 11762 3556 11886
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 3169 11387 3477 11396
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3160 8514 3188 9114
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3068 8486 3188 8514
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2976 6914 3004 8434
rect 3068 8430 3096 8486
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2884 6886 3004 6914
rect 3068 6914 3096 8366
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 3169 8123 3477 8132
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3068 6886 3188 6914
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2884 4146 2912 6886
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 5710 3004 6734
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6390 3096 6598
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3160 6100 3188 6886
rect 3068 6072 3188 6100
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2976 4010 3004 5646
rect 3068 4078 3096 6072
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 3528 3602 3556 11698
rect 3606 11656 3662 11665
rect 3606 11591 3608 11600
rect 3660 11591 3662 11600
rect 3608 11562 3660 11568
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3620 5234 3648 11018
rect 3712 8498 3740 12378
rect 3804 8838 3832 14742
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 3712 2650 3740 7822
rect 3804 6866 3832 8366
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3804 5370 3832 6802
rect 3896 6798 3924 17682
rect 3988 17542 4016 19722
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 18034 4108 19654
rect 4080 18006 4200 18034
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3974 17232 4030 17241
rect 3974 17167 3976 17176
rect 4028 17167 4030 17176
rect 3976 17138 4028 17144
rect 3988 16658 4016 17138
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 4080 16522 4108 17070
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14414 4016 14894
rect 4080 14618 4108 16458
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 13870 4016 14350
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3988 12646 4016 13806
rect 4080 13462 4108 14554
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 11830 4016 12582
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3988 10130 4016 11766
rect 4080 11354 4108 12786
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 4080 10010 4108 11290
rect 3988 9982 4108 10010
rect 3988 9178 4016 9982
rect 4172 9874 4200 18006
rect 4264 14618 4292 23530
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4356 11762 4384 23802
rect 4436 22228 4488 22234
rect 4436 22170 4488 22176
rect 4448 20602 4476 22170
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4448 13938 4476 19450
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4250 10976 4306 10985
rect 4250 10911 4306 10920
rect 4264 10062 4292 10911
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4172 9846 4292 9874
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3988 6662 4016 8978
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3804 4690 3832 5306
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3804 3602 3832 4626
rect 4080 4622 4108 9551
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3804 3058 3832 3538
rect 4172 3194 4200 9318
rect 4264 3534 4292 9846
rect 4448 6914 4476 12242
rect 4540 10690 4568 26522
rect 4632 25906 4660 27406
rect 4712 26512 4764 26518
rect 4712 26454 4764 26460
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 4724 23866 4752 26454
rect 4816 24750 4844 29038
rect 5000 27130 5028 29038
rect 4988 27124 5040 27130
rect 4988 27066 5040 27072
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 4908 26382 4936 26862
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 5092 26314 5120 29038
rect 5264 28960 5316 28966
rect 5264 28902 5316 28908
rect 5080 26308 5132 26314
rect 5080 26250 5132 26256
rect 5080 25832 5132 25838
rect 5080 25774 5132 25780
rect 5092 24954 5120 25774
rect 5172 25696 5224 25702
rect 5172 25638 5224 25644
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4804 24744 4856 24750
rect 4804 24686 4856 24692
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4724 15502 4752 23666
rect 4816 21962 4844 24686
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 4816 19378 4844 21898
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4724 11898 4752 14010
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4540 10662 4660 10690
rect 4632 10266 4660 10662
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4816 8634 4844 18226
rect 4908 13530 4936 24754
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5000 22030 5028 24142
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 5000 21554 5028 21966
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 5092 21146 5120 24890
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5184 20942 5212 25638
rect 5276 23730 5304 28902
rect 5724 28688 5776 28694
rect 5724 28630 5776 28636
rect 5388 28316 5696 28325
rect 5388 28314 5394 28316
rect 5450 28314 5474 28316
rect 5530 28314 5554 28316
rect 5610 28314 5634 28316
rect 5690 28314 5696 28316
rect 5450 28262 5452 28314
rect 5632 28262 5634 28314
rect 5388 28260 5394 28262
rect 5450 28260 5474 28262
rect 5530 28260 5554 28262
rect 5610 28260 5634 28262
rect 5690 28260 5696 28262
rect 5388 28251 5696 28260
rect 5388 27228 5696 27237
rect 5388 27226 5394 27228
rect 5450 27226 5474 27228
rect 5530 27226 5554 27228
rect 5610 27226 5634 27228
rect 5690 27226 5696 27228
rect 5450 27174 5452 27226
rect 5632 27174 5634 27226
rect 5388 27172 5394 27174
rect 5450 27172 5474 27174
rect 5530 27172 5554 27174
rect 5610 27172 5634 27174
rect 5690 27172 5696 27174
rect 5388 27163 5696 27172
rect 5736 27010 5764 28630
rect 5816 27532 5868 27538
rect 5816 27474 5868 27480
rect 5644 26994 5764 27010
rect 5632 26988 5764 26994
rect 5684 26982 5764 26988
rect 5632 26930 5684 26936
rect 5388 26140 5696 26149
rect 5388 26138 5394 26140
rect 5450 26138 5474 26140
rect 5530 26138 5554 26140
rect 5610 26138 5634 26140
rect 5690 26138 5696 26140
rect 5450 26086 5452 26138
rect 5632 26086 5634 26138
rect 5388 26084 5394 26086
rect 5450 26084 5474 26086
rect 5530 26084 5554 26086
rect 5610 26084 5634 26086
rect 5690 26084 5696 26086
rect 5388 26075 5696 26084
rect 5736 25430 5764 26982
rect 5828 26382 5856 27474
rect 5908 26784 5960 26790
rect 5908 26726 5960 26732
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 5828 25498 5856 26318
rect 5816 25492 5868 25498
rect 5816 25434 5868 25440
rect 5724 25424 5776 25430
rect 5724 25366 5776 25372
rect 5388 25052 5696 25061
rect 5388 25050 5394 25052
rect 5450 25050 5474 25052
rect 5530 25050 5554 25052
rect 5610 25050 5634 25052
rect 5690 25050 5696 25052
rect 5450 24998 5452 25050
rect 5632 24998 5634 25050
rect 5388 24996 5394 24998
rect 5450 24996 5474 24998
rect 5530 24996 5554 24998
rect 5610 24996 5634 24998
rect 5690 24996 5696 24998
rect 5388 24987 5696 24996
rect 5388 23964 5696 23973
rect 5388 23962 5394 23964
rect 5450 23962 5474 23964
rect 5530 23962 5554 23964
rect 5610 23962 5634 23964
rect 5690 23962 5696 23964
rect 5450 23910 5452 23962
rect 5632 23910 5634 23962
rect 5388 23908 5394 23910
rect 5450 23908 5474 23910
rect 5530 23908 5554 23910
rect 5610 23908 5634 23910
rect 5690 23908 5696 23910
rect 5388 23899 5696 23908
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5388 22876 5696 22885
rect 5388 22874 5394 22876
rect 5450 22874 5474 22876
rect 5530 22874 5554 22876
rect 5610 22874 5634 22876
rect 5690 22874 5696 22876
rect 5450 22822 5452 22874
rect 5632 22822 5634 22874
rect 5388 22820 5394 22822
rect 5450 22820 5474 22822
rect 5530 22820 5554 22822
rect 5610 22820 5634 22822
rect 5690 22820 5696 22822
rect 5388 22811 5696 22820
rect 5736 22778 5764 25366
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 5828 24342 5856 25230
rect 5816 24336 5868 24342
rect 5816 24278 5868 24284
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5736 22234 5764 22714
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5828 21962 5856 24074
rect 5920 23322 5948 26726
rect 6104 26450 6132 32234
rect 6196 30326 6224 32846
rect 6380 31346 6408 34138
rect 6472 33998 6500 34546
rect 6460 33992 6512 33998
rect 6460 33934 6512 33940
rect 6472 31414 6500 33934
rect 6932 32434 6960 34614
rect 7208 34066 7236 36110
rect 7300 35894 7328 36178
rect 9827 35932 10135 35941
rect 9827 35930 9833 35932
rect 9889 35930 9913 35932
rect 9969 35930 9993 35932
rect 10049 35930 10073 35932
rect 10129 35930 10135 35932
rect 7300 35866 7420 35894
rect 9889 35878 9891 35930
rect 10071 35878 10073 35930
rect 9827 35876 9833 35878
rect 9889 35876 9913 35878
rect 9969 35876 9993 35878
rect 10049 35876 10073 35878
rect 10129 35876 10135 35878
rect 9827 35867 10135 35876
rect 14266 35932 14574 35941
rect 14266 35930 14272 35932
rect 14328 35930 14352 35932
rect 14408 35930 14432 35932
rect 14488 35930 14512 35932
rect 14568 35930 14574 35932
rect 14328 35878 14330 35930
rect 14510 35878 14512 35930
rect 14266 35876 14272 35878
rect 14328 35876 14352 35878
rect 14408 35876 14432 35878
rect 14488 35876 14512 35878
rect 14568 35876 14574 35878
rect 14266 35867 14574 35876
rect 18705 35932 19013 35941
rect 18705 35930 18711 35932
rect 18767 35930 18791 35932
rect 18847 35930 18871 35932
rect 18927 35930 18951 35932
rect 19007 35930 19013 35932
rect 18767 35878 18769 35930
rect 18949 35878 18951 35930
rect 18705 35876 18711 35878
rect 18767 35876 18791 35878
rect 18847 35876 18871 35878
rect 18927 35876 18951 35878
rect 19007 35876 19013 35878
rect 18705 35867 19013 35876
rect 7288 34604 7340 34610
rect 7288 34546 7340 34552
rect 7196 34060 7248 34066
rect 7196 34002 7248 34008
rect 7208 33114 7236 34002
rect 7300 33998 7328 34546
rect 7392 34202 7420 35866
rect 7608 35388 7916 35397
rect 7608 35386 7614 35388
rect 7670 35386 7694 35388
rect 7750 35386 7774 35388
rect 7830 35386 7854 35388
rect 7910 35386 7916 35388
rect 7670 35334 7672 35386
rect 7852 35334 7854 35386
rect 7608 35332 7614 35334
rect 7670 35332 7694 35334
rect 7750 35332 7774 35334
rect 7830 35332 7854 35334
rect 7910 35332 7916 35334
rect 7608 35323 7916 35332
rect 12047 35388 12355 35397
rect 12047 35386 12053 35388
rect 12109 35386 12133 35388
rect 12189 35386 12213 35388
rect 12269 35386 12293 35388
rect 12349 35386 12355 35388
rect 12109 35334 12111 35386
rect 12291 35334 12293 35386
rect 12047 35332 12053 35334
rect 12109 35332 12133 35334
rect 12189 35332 12213 35334
rect 12269 35332 12293 35334
rect 12349 35332 12355 35334
rect 12047 35323 12355 35332
rect 16486 35388 16794 35397
rect 16486 35386 16492 35388
rect 16548 35386 16572 35388
rect 16628 35386 16652 35388
rect 16708 35386 16732 35388
rect 16788 35386 16794 35388
rect 16548 35334 16550 35386
rect 16730 35334 16732 35386
rect 16486 35332 16492 35334
rect 16548 35332 16572 35334
rect 16628 35332 16652 35334
rect 16708 35332 16732 35334
rect 16788 35332 16794 35334
rect 16486 35323 16794 35332
rect 9827 34844 10135 34853
rect 9827 34842 9833 34844
rect 9889 34842 9913 34844
rect 9969 34842 9993 34844
rect 10049 34842 10073 34844
rect 10129 34842 10135 34844
rect 9889 34790 9891 34842
rect 10071 34790 10073 34842
rect 9827 34788 9833 34790
rect 9889 34788 9913 34790
rect 9969 34788 9993 34790
rect 10049 34788 10073 34790
rect 10129 34788 10135 34790
rect 9827 34779 10135 34788
rect 14266 34844 14574 34853
rect 14266 34842 14272 34844
rect 14328 34842 14352 34844
rect 14408 34842 14432 34844
rect 14488 34842 14512 34844
rect 14568 34842 14574 34844
rect 14328 34790 14330 34842
rect 14510 34790 14512 34842
rect 14266 34788 14272 34790
rect 14328 34788 14352 34790
rect 14408 34788 14432 34790
rect 14488 34788 14512 34790
rect 14568 34788 14574 34790
rect 14266 34779 14574 34788
rect 18705 34844 19013 34853
rect 18705 34842 18711 34844
rect 18767 34842 18791 34844
rect 18847 34842 18871 34844
rect 18927 34842 18951 34844
rect 19007 34842 19013 34844
rect 18767 34790 18769 34842
rect 18949 34790 18951 34842
rect 18705 34788 18711 34790
rect 18767 34788 18791 34790
rect 18847 34788 18871 34790
rect 18927 34788 18951 34790
rect 19007 34788 19013 34790
rect 18705 34779 19013 34788
rect 7608 34300 7916 34309
rect 7608 34298 7614 34300
rect 7670 34298 7694 34300
rect 7750 34298 7774 34300
rect 7830 34298 7854 34300
rect 7910 34298 7916 34300
rect 7670 34246 7672 34298
rect 7852 34246 7854 34298
rect 7608 34244 7614 34246
rect 7670 34244 7694 34246
rect 7750 34244 7774 34246
rect 7830 34244 7854 34246
rect 7910 34244 7916 34246
rect 7608 34235 7916 34244
rect 12047 34300 12355 34309
rect 12047 34298 12053 34300
rect 12109 34298 12133 34300
rect 12189 34298 12213 34300
rect 12269 34298 12293 34300
rect 12349 34298 12355 34300
rect 12109 34246 12111 34298
rect 12291 34246 12293 34298
rect 12047 34244 12053 34246
rect 12109 34244 12133 34246
rect 12189 34244 12213 34246
rect 12269 34244 12293 34246
rect 12349 34244 12355 34246
rect 12047 34235 12355 34244
rect 16486 34300 16794 34309
rect 16486 34298 16492 34300
rect 16548 34298 16572 34300
rect 16628 34298 16652 34300
rect 16708 34298 16732 34300
rect 16788 34298 16794 34300
rect 16548 34246 16550 34298
rect 16730 34246 16732 34298
rect 16486 34244 16492 34246
rect 16548 34244 16572 34246
rect 16628 34244 16652 34246
rect 16708 34244 16732 34246
rect 16788 34244 16794 34246
rect 16486 34235 16794 34244
rect 7380 34196 7432 34202
rect 7380 34138 7432 34144
rect 7288 33992 7340 33998
rect 7288 33934 7340 33940
rect 7196 33108 7248 33114
rect 7196 33050 7248 33056
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 6828 32428 6880 32434
rect 6828 32370 6880 32376
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6460 31408 6512 31414
rect 6460 31350 6512 31356
rect 6368 31340 6420 31346
rect 6368 31282 6420 31288
rect 6472 30870 6500 31350
rect 6460 30864 6512 30870
rect 6460 30806 6512 30812
rect 6368 30728 6420 30734
rect 6368 30670 6420 30676
rect 6184 30320 6236 30326
rect 6184 30262 6236 30268
rect 6196 29646 6224 30262
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6196 27062 6224 29582
rect 6380 28506 6408 30670
rect 6552 30660 6604 30666
rect 6552 30602 6604 30608
rect 6460 29028 6512 29034
rect 6460 28970 6512 28976
rect 6472 28626 6500 28970
rect 6460 28620 6512 28626
rect 6460 28562 6512 28568
rect 6564 28558 6592 30602
rect 6656 29170 6684 32166
rect 6840 31754 6868 32370
rect 7116 31754 7144 32846
rect 7300 31754 7328 33934
rect 6748 31726 6868 31754
rect 7024 31726 7144 31754
rect 7208 31726 7328 31754
rect 6748 30394 6776 31726
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 6736 30388 6788 30394
rect 6736 30330 6788 30336
rect 6748 29646 6776 30330
rect 6840 30054 6868 31282
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6840 29170 6868 29990
rect 6932 29306 6960 30534
rect 7024 30258 7052 31726
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 7012 30252 7064 30258
rect 7012 30194 7064 30200
rect 7024 29782 7052 30194
rect 7012 29776 7064 29782
rect 7012 29718 7064 29724
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 6920 29300 6972 29306
rect 6920 29242 6972 29248
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6736 29096 6788 29102
rect 6736 29038 6788 29044
rect 6748 28558 6776 29038
rect 6840 28626 6868 29106
rect 6828 28620 6880 28626
rect 6828 28562 6880 28568
rect 6552 28552 6604 28558
rect 6380 28478 6500 28506
rect 6552 28494 6604 28500
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 6276 28416 6328 28422
rect 6276 28358 6328 28364
rect 6184 27056 6236 27062
rect 6184 26998 6236 27004
rect 6288 26518 6316 28358
rect 6472 28082 6500 28478
rect 6460 28076 6512 28082
rect 6460 28018 6512 28024
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6276 26512 6328 26518
rect 6276 26454 6328 26460
rect 6092 26444 6144 26450
rect 6092 26386 6144 26392
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 6182 26344 6238 26353
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5724 21956 5776 21962
rect 5724 21898 5776 21904
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5736 21842 5764 21898
rect 5276 21690 5304 21830
rect 5736 21814 5856 21842
rect 5388 21788 5696 21797
rect 5388 21786 5394 21788
rect 5450 21786 5474 21788
rect 5530 21786 5554 21788
rect 5610 21786 5634 21788
rect 5690 21786 5696 21788
rect 5450 21734 5452 21786
rect 5632 21734 5634 21786
rect 5388 21732 5394 21734
rect 5450 21732 5474 21734
rect 5530 21732 5554 21734
rect 5610 21732 5634 21734
rect 5690 21732 5696 21734
rect 5388 21723 5696 21732
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5828 21554 5856 21814
rect 5920 21622 5948 23258
rect 6012 23254 6040 26318
rect 6182 26279 6184 26288
rect 6236 26279 6238 26288
rect 6184 26250 6236 26256
rect 6380 25226 6408 26930
rect 6472 26382 6500 28018
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6276 24404 6328 24410
rect 6276 24346 6328 24352
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6000 23248 6052 23254
rect 6000 23190 6052 23196
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6012 22778 6040 23054
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5908 21616 5960 21622
rect 5908 21558 5960 21564
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 5276 20466 5304 21490
rect 5388 20700 5696 20709
rect 5388 20698 5394 20700
rect 5450 20698 5474 20700
rect 5530 20698 5554 20700
rect 5610 20698 5634 20700
rect 5690 20698 5696 20700
rect 5450 20646 5452 20698
rect 5632 20646 5634 20698
rect 5388 20644 5394 20646
rect 5450 20644 5474 20646
rect 5530 20644 5554 20646
rect 5610 20644 5634 20646
rect 5690 20644 5696 20646
rect 5388 20635 5696 20644
rect 5736 20534 5764 21490
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 5828 20466 5856 21490
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 5920 20874 5948 21422
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4448 6886 4660 6914
rect 4632 6458 4660 6886
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4802 5536 4858 5545
rect 4802 5471 4858 5480
rect 4816 4622 4844 5471
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4908 4146 4936 6054
rect 5000 5098 5028 16458
rect 5276 16250 5304 20402
rect 5388 19612 5696 19621
rect 5388 19610 5394 19612
rect 5450 19610 5474 19612
rect 5530 19610 5554 19612
rect 5610 19610 5634 19612
rect 5690 19610 5696 19612
rect 5450 19558 5452 19610
rect 5632 19558 5634 19610
rect 5388 19556 5394 19558
rect 5450 19556 5474 19558
rect 5530 19556 5554 19558
rect 5610 19556 5634 19558
rect 5690 19556 5696 19558
rect 5388 19547 5696 19556
rect 5724 19440 5776 19446
rect 5724 19382 5776 19388
rect 5388 18524 5696 18533
rect 5388 18522 5394 18524
rect 5450 18522 5474 18524
rect 5530 18522 5554 18524
rect 5610 18522 5634 18524
rect 5690 18522 5696 18524
rect 5450 18470 5452 18522
rect 5632 18470 5634 18522
rect 5388 18468 5394 18470
rect 5450 18468 5474 18470
rect 5530 18468 5554 18470
rect 5610 18468 5634 18470
rect 5690 18468 5696 18470
rect 5388 18459 5696 18468
rect 5388 17436 5696 17445
rect 5388 17434 5394 17436
rect 5450 17434 5474 17436
rect 5530 17434 5554 17436
rect 5610 17434 5634 17436
rect 5690 17434 5696 17436
rect 5450 17382 5452 17434
rect 5632 17382 5634 17434
rect 5388 17380 5394 17382
rect 5450 17380 5474 17382
rect 5530 17380 5554 17382
rect 5610 17380 5634 17382
rect 5690 17380 5696 17382
rect 5388 17371 5696 17380
rect 5388 16348 5696 16357
rect 5388 16346 5394 16348
rect 5450 16346 5474 16348
rect 5530 16346 5554 16348
rect 5610 16346 5634 16348
rect 5690 16346 5696 16348
rect 5450 16294 5452 16346
rect 5632 16294 5634 16346
rect 5388 16292 5394 16294
rect 5450 16292 5474 16294
rect 5530 16292 5554 16294
rect 5610 16292 5634 16294
rect 5690 16292 5696 16294
rect 5388 16283 5696 16292
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3804 2514 3832 2994
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 1952 2372 2004 2378
rect 1952 2314 2004 2320
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 5000 800 5028 3470
rect 5092 2446 5120 15302
rect 5388 15260 5696 15269
rect 5388 15258 5394 15260
rect 5450 15258 5474 15260
rect 5530 15258 5554 15260
rect 5610 15258 5634 15260
rect 5690 15258 5696 15260
rect 5450 15206 5452 15258
rect 5632 15206 5634 15258
rect 5388 15204 5394 15206
rect 5450 15204 5474 15206
rect 5530 15204 5554 15206
rect 5610 15204 5634 15206
rect 5690 15204 5696 15206
rect 5388 15195 5696 15204
rect 5736 15162 5764 19382
rect 5920 18766 5948 20810
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5828 15450 5856 16526
rect 5908 15496 5960 15502
rect 5828 15444 5908 15450
rect 5828 15438 5960 15444
rect 5828 15422 5948 15438
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5828 14958 5856 15422
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5276 14074 5304 14282
rect 5388 14172 5696 14181
rect 5388 14170 5394 14172
rect 5450 14170 5474 14172
rect 5530 14170 5554 14172
rect 5610 14170 5634 14172
rect 5690 14170 5696 14172
rect 5450 14118 5452 14170
rect 5632 14118 5634 14170
rect 5388 14116 5394 14118
rect 5450 14116 5474 14118
rect 5530 14116 5554 14118
rect 5610 14116 5634 14118
rect 5690 14116 5696 14118
rect 5388 14107 5696 14116
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5170 13832 5226 13841
rect 5170 13767 5226 13776
rect 5184 6798 5212 13767
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5276 12850 5304 13194
rect 5388 13084 5696 13093
rect 5388 13082 5394 13084
rect 5450 13082 5474 13084
rect 5530 13082 5554 13084
rect 5610 13082 5634 13084
rect 5690 13082 5696 13084
rect 5450 13030 5452 13082
rect 5632 13030 5634 13082
rect 5388 13028 5394 13030
rect 5450 13028 5474 13030
rect 5530 13028 5554 13030
rect 5610 13028 5634 13030
rect 5690 13028 5696 13030
rect 5388 13019 5696 13028
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5276 10198 5304 12786
rect 5388 11996 5696 12005
rect 5388 11994 5394 11996
rect 5450 11994 5474 11996
rect 5530 11994 5554 11996
rect 5610 11994 5634 11996
rect 5690 11994 5696 11996
rect 5450 11942 5452 11994
rect 5632 11942 5634 11994
rect 5388 11940 5394 11942
rect 5450 11940 5474 11942
rect 5530 11940 5554 11942
rect 5610 11940 5634 11942
rect 5690 11940 5696 11942
rect 5388 11931 5696 11940
rect 5736 11762 5764 14554
rect 5828 14414 5856 14894
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5920 14074 5948 15098
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6012 12434 6040 22578
rect 6104 22030 6132 24142
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 6196 22098 6224 23122
rect 6184 22092 6236 22098
rect 6288 22094 6316 24346
rect 6380 23866 6408 25162
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 6380 22710 6408 23802
rect 6368 22704 6420 22710
rect 6368 22646 6420 22652
rect 6288 22066 6408 22094
rect 6184 22034 6236 22040
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6184 21956 6236 21962
rect 6184 21898 6236 21904
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6104 21690 6132 21830
rect 6092 21684 6144 21690
rect 6092 21626 6144 21632
rect 6092 20528 6144 20534
rect 6092 20470 6144 20476
rect 5920 12406 6040 12434
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5388 10908 5696 10917
rect 5388 10906 5394 10908
rect 5450 10906 5474 10908
rect 5530 10906 5554 10908
rect 5610 10906 5634 10908
rect 5690 10906 5696 10908
rect 5450 10854 5452 10906
rect 5632 10854 5634 10906
rect 5388 10852 5394 10854
rect 5450 10852 5474 10854
rect 5530 10852 5554 10854
rect 5610 10852 5634 10854
rect 5690 10852 5696 10854
rect 5388 10843 5696 10852
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5276 5710 5304 10134
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5388 9820 5696 9829
rect 5388 9818 5394 9820
rect 5450 9818 5474 9820
rect 5530 9818 5554 9820
rect 5610 9818 5634 9820
rect 5690 9818 5696 9820
rect 5450 9766 5452 9818
rect 5632 9766 5634 9818
rect 5388 9764 5394 9766
rect 5450 9764 5474 9766
rect 5530 9764 5554 9766
rect 5610 9764 5634 9766
rect 5690 9764 5696 9766
rect 5388 9755 5696 9764
rect 5388 8732 5696 8741
rect 5388 8730 5394 8732
rect 5450 8730 5474 8732
rect 5530 8730 5554 8732
rect 5610 8730 5634 8732
rect 5690 8730 5696 8732
rect 5450 8678 5452 8730
rect 5632 8678 5634 8730
rect 5388 8676 5394 8678
rect 5450 8676 5474 8678
rect 5530 8676 5554 8678
rect 5610 8676 5634 8678
rect 5690 8676 5696 8678
rect 5388 8667 5696 8676
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5276 5302 5304 5646
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 5828 3534 5856 9930
rect 5920 6914 5948 12406
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 11218 6040 12242
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10674 6040 11154
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5920 6886 6040 6914
rect 6012 4486 6040 6886
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6104 4078 6132 20470
rect 6196 16250 6224 21898
rect 6380 21894 6408 22066
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6288 16114 6316 20334
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6196 15502 6224 15982
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6196 14958 6224 15438
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6196 14414 6224 14894
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13870 6224 14350
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6288 7002 6316 14962
rect 6380 10810 6408 20402
rect 6472 18970 6500 26318
rect 6564 24206 6592 28494
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6656 24750 6684 27270
rect 6840 27062 6868 27338
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 6736 26852 6788 26858
rect 6736 26794 6788 26800
rect 6748 25158 6776 26794
rect 6840 25974 6868 26998
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6828 25968 6880 25974
rect 6828 25910 6880 25916
rect 6932 25838 6960 26862
rect 7024 26042 7052 29582
rect 7116 29170 7144 31282
rect 7208 30666 7236 31726
rect 7288 31272 7340 31278
rect 7288 31214 7340 31220
rect 7196 30660 7248 30666
rect 7196 30602 7248 30608
rect 7196 30184 7248 30190
rect 7196 30126 7248 30132
rect 7104 29164 7156 29170
rect 7104 29106 7156 29112
rect 7012 26036 7064 26042
rect 7012 25978 7064 25984
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 6828 25220 6880 25226
rect 6828 25162 6880 25168
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6644 24744 6696 24750
rect 6644 24686 6696 24692
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6564 23050 6592 23598
rect 6552 23044 6604 23050
rect 6552 22986 6604 22992
rect 6564 20398 6592 22986
rect 6656 22642 6684 24686
rect 6748 24410 6776 25094
rect 6840 24886 6868 25162
rect 6828 24880 6880 24886
rect 6828 24822 6880 24828
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6840 22778 6868 24822
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6826 20768 6882 20777
rect 6826 20703 6882 20712
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6472 14414 6500 15914
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6472 13190 6500 13806
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6472 12782 6500 13126
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6472 12306 6500 12718
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6472 4622 6500 11698
rect 6564 8566 6592 20198
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 9654 6684 18634
rect 6840 15094 6868 20703
rect 6932 18698 6960 25774
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 7024 24274 7052 25298
rect 7116 24682 7144 29106
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 7010 24168 7066 24177
rect 7010 24103 7066 24112
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6564 5914 6592 6258
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6564 5234 6592 5850
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6564 4826 6592 5170
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6564 4146 6592 4762
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6288 3602 6316 4082
rect 6748 3738 6776 12038
rect 6826 6624 6882 6633
rect 6826 6559 6882 6568
rect 6840 6322 6868 6559
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6840 4146 6868 5850
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 7024 3602 7052 24103
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7116 22982 7144 23666
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7116 22234 7144 22578
rect 7208 22234 7236 30126
rect 7300 28558 7328 31214
rect 7392 30122 7420 34138
rect 8668 34128 8720 34134
rect 8668 34070 8720 34076
rect 7608 33212 7916 33221
rect 7608 33210 7614 33212
rect 7670 33210 7694 33212
rect 7750 33210 7774 33212
rect 7830 33210 7854 33212
rect 7910 33210 7916 33212
rect 7670 33158 7672 33210
rect 7852 33158 7854 33210
rect 7608 33156 7614 33158
rect 7670 33156 7694 33158
rect 7750 33156 7774 33158
rect 7830 33156 7854 33158
rect 7910 33156 7916 33158
rect 7608 33147 7916 33156
rect 7932 32768 7984 32774
rect 7932 32710 7984 32716
rect 7608 32124 7916 32133
rect 7608 32122 7614 32124
rect 7670 32122 7694 32124
rect 7750 32122 7774 32124
rect 7830 32122 7854 32124
rect 7910 32122 7916 32124
rect 7670 32070 7672 32122
rect 7852 32070 7854 32122
rect 7608 32068 7614 32070
rect 7670 32068 7694 32070
rect 7750 32068 7774 32070
rect 7830 32068 7854 32070
rect 7910 32068 7916 32070
rect 7608 32059 7916 32068
rect 7608 31036 7916 31045
rect 7608 31034 7614 31036
rect 7670 31034 7694 31036
rect 7750 31034 7774 31036
rect 7830 31034 7854 31036
rect 7910 31034 7916 31036
rect 7670 30982 7672 31034
rect 7852 30982 7854 31034
rect 7608 30980 7614 30982
rect 7670 30980 7694 30982
rect 7750 30980 7774 30982
rect 7830 30980 7854 30982
rect 7910 30980 7916 30982
rect 7608 30971 7916 30980
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7380 30116 7432 30122
rect 7380 30058 7432 30064
rect 7484 29850 7512 30670
rect 7564 30660 7616 30666
rect 7564 30602 7616 30608
rect 7576 30394 7604 30602
rect 7564 30388 7616 30394
rect 7564 30330 7616 30336
rect 7944 30258 7972 32710
rect 8024 30592 8076 30598
rect 8024 30534 8076 30540
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 8036 30138 8064 30534
rect 7944 30110 8064 30138
rect 7608 29948 7916 29957
rect 7608 29946 7614 29948
rect 7670 29946 7694 29948
rect 7750 29946 7774 29948
rect 7830 29946 7854 29948
rect 7910 29946 7916 29948
rect 7670 29894 7672 29946
rect 7852 29894 7854 29946
rect 7608 29892 7614 29894
rect 7670 29892 7694 29894
rect 7750 29892 7774 29894
rect 7830 29892 7854 29894
rect 7910 29892 7916 29894
rect 7608 29883 7916 29892
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7300 28422 7328 28494
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7300 26382 7328 28358
rect 7392 26926 7420 29582
rect 7484 29306 7512 29786
rect 7472 29300 7524 29306
rect 7472 29242 7524 29248
rect 7472 29164 7524 29170
rect 7472 29106 7524 29112
rect 7484 28558 7512 29106
rect 7608 28860 7916 28869
rect 7608 28858 7614 28860
rect 7670 28858 7694 28860
rect 7750 28858 7774 28860
rect 7830 28858 7854 28860
rect 7910 28858 7916 28860
rect 7670 28806 7672 28858
rect 7852 28806 7854 28858
rect 7608 28804 7614 28806
rect 7670 28804 7694 28806
rect 7750 28804 7774 28806
rect 7830 28804 7854 28806
rect 7910 28804 7916 28806
rect 7608 28795 7916 28804
rect 7944 28558 7972 30110
rect 8116 30048 8168 30054
rect 8116 29990 8168 29996
rect 8024 29164 8076 29170
rect 8024 29106 8076 29112
rect 7472 28552 7524 28558
rect 7472 28494 7524 28500
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7484 27169 7512 28494
rect 7608 27772 7916 27781
rect 7608 27770 7614 27772
rect 7670 27770 7694 27772
rect 7750 27770 7774 27772
rect 7830 27770 7854 27772
rect 7910 27770 7916 27772
rect 7670 27718 7672 27770
rect 7852 27718 7854 27770
rect 7608 27716 7614 27718
rect 7670 27716 7694 27718
rect 7750 27716 7774 27718
rect 7830 27716 7854 27718
rect 7910 27716 7916 27718
rect 7608 27707 7916 27716
rect 7470 27160 7526 27169
rect 7470 27095 7526 27104
rect 7472 27056 7524 27062
rect 7472 26998 7524 27004
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7300 24206 7328 26318
rect 7392 25838 7420 26862
rect 7484 25906 7512 26998
rect 7608 26684 7916 26693
rect 7608 26682 7614 26684
rect 7670 26682 7694 26684
rect 7750 26682 7774 26684
rect 7830 26682 7854 26684
rect 7910 26682 7916 26684
rect 7670 26630 7672 26682
rect 7852 26630 7854 26682
rect 7608 26628 7614 26630
rect 7670 26628 7694 26630
rect 7750 26628 7774 26630
rect 7830 26628 7854 26630
rect 7910 26628 7916 26630
rect 7608 26619 7916 26628
rect 7944 26314 7972 28494
rect 8036 28014 8064 29106
rect 8128 29073 8156 29990
rect 8208 29776 8260 29782
rect 8208 29718 8260 29724
rect 8114 29064 8170 29073
rect 8114 28999 8170 29008
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 7932 26308 7984 26314
rect 7932 26250 7984 26256
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 7392 24698 7420 25774
rect 7608 25596 7916 25605
rect 7608 25594 7614 25596
rect 7670 25594 7694 25596
rect 7750 25594 7774 25596
rect 7830 25594 7854 25596
rect 7910 25594 7916 25596
rect 7670 25542 7672 25594
rect 7852 25542 7854 25594
rect 7608 25540 7614 25542
rect 7670 25540 7694 25542
rect 7750 25540 7774 25542
rect 7830 25540 7854 25542
rect 7910 25540 7916 25542
rect 7608 25531 7916 25540
rect 7840 25288 7892 25294
rect 7838 25256 7840 25265
rect 7892 25256 7894 25265
rect 7838 25191 7894 25200
rect 8036 24818 8064 27950
rect 8220 26246 8248 29718
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 8208 26240 8260 26246
rect 8208 26182 8260 26188
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 7932 24744 7984 24750
rect 7392 24670 7604 24698
rect 7932 24686 7984 24692
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 7196 22228 7248 22234
rect 7196 22170 7248 22176
rect 7116 22030 7144 22170
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 12986 7144 16934
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7208 7546 7236 20742
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7116 6390 7144 6666
rect 7300 6458 7328 22714
rect 7392 22710 7420 24670
rect 7576 24614 7604 24670
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7484 23730 7512 24550
rect 7608 24508 7916 24517
rect 7608 24506 7614 24508
rect 7670 24506 7694 24508
rect 7750 24506 7774 24508
rect 7830 24506 7854 24508
rect 7910 24506 7916 24508
rect 7670 24454 7672 24506
rect 7852 24454 7854 24506
rect 7608 24452 7614 24454
rect 7670 24452 7694 24454
rect 7750 24452 7774 24454
rect 7830 24452 7854 24454
rect 7910 24452 7916 24454
rect 7608 24443 7916 24452
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7852 24206 7880 24346
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7944 23730 7972 24686
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7484 22642 7512 23666
rect 7608 23420 7916 23429
rect 7608 23418 7614 23420
rect 7670 23418 7694 23420
rect 7750 23418 7774 23420
rect 7830 23418 7854 23420
rect 7910 23418 7916 23420
rect 7670 23366 7672 23418
rect 7852 23366 7854 23418
rect 7608 23364 7614 23366
rect 7670 23364 7694 23366
rect 7750 23364 7774 23366
rect 7830 23364 7854 23366
rect 7910 23364 7916 23366
rect 7608 23355 7916 23364
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7484 22522 7512 22578
rect 7944 22522 7972 23666
rect 7392 22494 7512 22522
rect 7852 22494 7972 22522
rect 7392 21962 7420 22494
rect 7852 22438 7880 22494
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7392 4554 7420 21898
rect 7484 20942 7512 22374
rect 7608 22332 7916 22341
rect 7608 22330 7614 22332
rect 7670 22330 7694 22332
rect 7750 22330 7774 22332
rect 7830 22330 7854 22332
rect 7910 22330 7916 22332
rect 7670 22278 7672 22330
rect 7852 22278 7854 22330
rect 7608 22276 7614 22278
rect 7670 22276 7694 22278
rect 7750 22276 7774 22278
rect 7830 22276 7854 22278
rect 7910 22276 7916 22278
rect 7608 22267 7916 22276
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7852 21622 7880 21898
rect 7840 21616 7892 21622
rect 7840 21558 7892 21564
rect 7608 21244 7916 21253
rect 7608 21242 7614 21244
rect 7670 21242 7694 21244
rect 7750 21242 7774 21244
rect 7830 21242 7854 21244
rect 7910 21242 7916 21244
rect 7670 21190 7672 21242
rect 7852 21190 7854 21242
rect 7608 21188 7614 21190
rect 7670 21188 7694 21190
rect 7750 21188 7774 21190
rect 7830 21188 7854 21190
rect 7910 21188 7916 21190
rect 7608 21179 7916 21188
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7484 20806 7512 20878
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7608 20156 7916 20165
rect 7608 20154 7614 20156
rect 7670 20154 7694 20156
rect 7750 20154 7774 20156
rect 7830 20154 7854 20156
rect 7910 20154 7916 20156
rect 7670 20102 7672 20154
rect 7852 20102 7854 20154
rect 7608 20100 7614 20102
rect 7670 20100 7694 20102
rect 7750 20100 7774 20102
rect 7830 20100 7854 20102
rect 7910 20100 7916 20102
rect 7608 20091 7916 20100
rect 7608 19068 7916 19077
rect 7608 19066 7614 19068
rect 7670 19066 7694 19068
rect 7750 19066 7774 19068
rect 7830 19066 7854 19068
rect 7910 19066 7916 19068
rect 7670 19014 7672 19066
rect 7852 19014 7854 19066
rect 7608 19012 7614 19014
rect 7670 19012 7694 19014
rect 7750 19012 7774 19014
rect 7830 19012 7854 19014
rect 7910 19012 7916 19014
rect 7608 19003 7916 19012
rect 7608 17980 7916 17989
rect 7608 17978 7614 17980
rect 7670 17978 7694 17980
rect 7750 17978 7774 17980
rect 7830 17978 7854 17980
rect 7910 17978 7916 17980
rect 7670 17926 7672 17978
rect 7852 17926 7854 17978
rect 7608 17924 7614 17926
rect 7670 17924 7694 17926
rect 7750 17924 7774 17926
rect 7830 17924 7854 17926
rect 7910 17924 7916 17926
rect 7608 17915 7916 17924
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7484 15706 7512 16730
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7944 15026 7972 22374
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 7608 13628 7916 13637
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 8036 9518 8064 24754
rect 8128 22778 8156 25434
rect 8312 25226 8340 26794
rect 8484 26784 8536 26790
rect 8484 26726 8536 26732
rect 8392 26240 8444 26246
rect 8392 26182 8444 26188
rect 8300 25220 8352 25226
rect 8300 25162 8352 25168
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 8128 15162 8156 22170
rect 8220 21962 8248 25094
rect 8312 23322 8340 25162
rect 8404 24886 8432 26182
rect 8392 24880 8444 24886
rect 8392 24822 8444 24828
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 8312 22778 8340 22918
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8220 21146 8248 21490
rect 8312 21350 8340 22578
rect 8392 21412 8444 21418
rect 8392 21354 8444 21360
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 8128 5370 8156 14962
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 7410 8248 9454
rect 8404 7478 8432 21354
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 6730 8248 7346
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8496 5914 8524 26726
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8588 5302 8616 26250
rect 8680 12918 8708 34070
rect 9827 33756 10135 33765
rect 9827 33754 9833 33756
rect 9889 33754 9913 33756
rect 9969 33754 9993 33756
rect 10049 33754 10073 33756
rect 10129 33754 10135 33756
rect 9889 33702 9891 33754
rect 10071 33702 10073 33754
rect 9827 33700 9833 33702
rect 9889 33700 9913 33702
rect 9969 33700 9993 33702
rect 10049 33700 10073 33702
rect 10129 33700 10135 33702
rect 9827 33691 10135 33700
rect 14266 33756 14574 33765
rect 14266 33754 14272 33756
rect 14328 33754 14352 33756
rect 14408 33754 14432 33756
rect 14488 33754 14512 33756
rect 14568 33754 14574 33756
rect 14328 33702 14330 33754
rect 14510 33702 14512 33754
rect 14266 33700 14272 33702
rect 14328 33700 14352 33702
rect 14408 33700 14432 33702
rect 14488 33700 14512 33702
rect 14568 33700 14574 33702
rect 14266 33691 14574 33700
rect 18705 33756 19013 33765
rect 18705 33754 18711 33756
rect 18767 33754 18791 33756
rect 18847 33754 18871 33756
rect 18927 33754 18951 33756
rect 19007 33754 19013 33756
rect 18767 33702 18769 33754
rect 18949 33702 18951 33754
rect 18705 33700 18711 33702
rect 18767 33700 18791 33702
rect 18847 33700 18871 33702
rect 18927 33700 18951 33702
rect 19007 33700 19013 33702
rect 18705 33691 19013 33700
rect 12047 33212 12355 33221
rect 12047 33210 12053 33212
rect 12109 33210 12133 33212
rect 12189 33210 12213 33212
rect 12269 33210 12293 33212
rect 12349 33210 12355 33212
rect 12109 33158 12111 33210
rect 12291 33158 12293 33210
rect 12047 33156 12053 33158
rect 12109 33156 12133 33158
rect 12189 33156 12213 33158
rect 12269 33156 12293 33158
rect 12349 33156 12355 33158
rect 12047 33147 12355 33156
rect 16486 33212 16794 33221
rect 16486 33210 16492 33212
rect 16548 33210 16572 33212
rect 16628 33210 16652 33212
rect 16708 33210 16732 33212
rect 16788 33210 16794 33212
rect 16548 33158 16550 33210
rect 16730 33158 16732 33210
rect 16486 33156 16492 33158
rect 16548 33156 16572 33158
rect 16628 33156 16652 33158
rect 16708 33156 16732 33158
rect 16788 33156 16794 33158
rect 16486 33147 16794 33156
rect 9827 32668 10135 32677
rect 9827 32666 9833 32668
rect 9889 32666 9913 32668
rect 9969 32666 9993 32668
rect 10049 32666 10073 32668
rect 10129 32666 10135 32668
rect 9889 32614 9891 32666
rect 10071 32614 10073 32666
rect 9827 32612 9833 32614
rect 9889 32612 9913 32614
rect 9969 32612 9993 32614
rect 10049 32612 10073 32614
rect 10129 32612 10135 32614
rect 9827 32603 10135 32612
rect 14266 32668 14574 32677
rect 14266 32666 14272 32668
rect 14328 32666 14352 32668
rect 14408 32666 14432 32668
rect 14488 32666 14512 32668
rect 14568 32666 14574 32668
rect 14328 32614 14330 32666
rect 14510 32614 14512 32666
rect 14266 32612 14272 32614
rect 14328 32612 14352 32614
rect 14408 32612 14432 32614
rect 14488 32612 14512 32614
rect 14568 32612 14574 32614
rect 14266 32603 14574 32612
rect 18705 32668 19013 32677
rect 18705 32666 18711 32668
rect 18767 32666 18791 32668
rect 18847 32666 18871 32668
rect 18927 32666 18951 32668
rect 19007 32666 19013 32668
rect 18767 32614 18769 32666
rect 18949 32614 18951 32666
rect 18705 32612 18711 32614
rect 18767 32612 18791 32614
rect 18847 32612 18871 32614
rect 18927 32612 18951 32614
rect 19007 32612 19013 32614
rect 18705 32603 19013 32612
rect 12047 32124 12355 32133
rect 12047 32122 12053 32124
rect 12109 32122 12133 32124
rect 12189 32122 12213 32124
rect 12269 32122 12293 32124
rect 12349 32122 12355 32124
rect 12109 32070 12111 32122
rect 12291 32070 12293 32122
rect 12047 32068 12053 32070
rect 12109 32068 12133 32070
rect 12189 32068 12213 32070
rect 12269 32068 12293 32070
rect 12349 32068 12355 32070
rect 12047 32059 12355 32068
rect 16486 32124 16794 32133
rect 16486 32122 16492 32124
rect 16548 32122 16572 32124
rect 16628 32122 16652 32124
rect 16708 32122 16732 32124
rect 16788 32122 16794 32124
rect 16548 32070 16550 32122
rect 16730 32070 16732 32122
rect 16486 32068 16492 32070
rect 16548 32068 16572 32070
rect 16628 32068 16652 32070
rect 16708 32068 16732 32070
rect 16788 32068 16794 32070
rect 16486 32059 16794 32068
rect 9827 31580 10135 31589
rect 9827 31578 9833 31580
rect 9889 31578 9913 31580
rect 9969 31578 9993 31580
rect 10049 31578 10073 31580
rect 10129 31578 10135 31580
rect 9889 31526 9891 31578
rect 10071 31526 10073 31578
rect 9827 31524 9833 31526
rect 9889 31524 9913 31526
rect 9969 31524 9993 31526
rect 10049 31524 10073 31526
rect 10129 31524 10135 31526
rect 9827 31515 10135 31524
rect 14266 31580 14574 31589
rect 14266 31578 14272 31580
rect 14328 31578 14352 31580
rect 14408 31578 14432 31580
rect 14488 31578 14512 31580
rect 14568 31578 14574 31580
rect 14328 31526 14330 31578
rect 14510 31526 14512 31578
rect 14266 31524 14272 31526
rect 14328 31524 14352 31526
rect 14408 31524 14432 31526
rect 14488 31524 14512 31526
rect 14568 31524 14574 31526
rect 14266 31515 14574 31524
rect 18705 31580 19013 31589
rect 18705 31578 18711 31580
rect 18767 31578 18791 31580
rect 18847 31578 18871 31580
rect 18927 31578 18951 31580
rect 19007 31578 19013 31580
rect 18767 31526 18769 31578
rect 18949 31526 18951 31578
rect 18705 31524 18711 31526
rect 18767 31524 18791 31526
rect 18847 31524 18871 31526
rect 18927 31524 18951 31526
rect 19007 31524 19013 31526
rect 18705 31515 19013 31524
rect 8852 31136 8904 31142
rect 8852 31078 8904 31084
rect 8760 26512 8812 26518
rect 8760 26454 8812 26460
rect 8772 13938 8800 26454
rect 8864 15366 8892 31078
rect 12047 31036 12355 31045
rect 12047 31034 12053 31036
rect 12109 31034 12133 31036
rect 12189 31034 12213 31036
rect 12269 31034 12293 31036
rect 12349 31034 12355 31036
rect 12109 30982 12111 31034
rect 12291 30982 12293 31034
rect 12047 30980 12053 30982
rect 12109 30980 12133 30982
rect 12189 30980 12213 30982
rect 12269 30980 12293 30982
rect 12349 30980 12355 30982
rect 12047 30971 12355 30980
rect 16486 31036 16794 31045
rect 16486 31034 16492 31036
rect 16548 31034 16572 31036
rect 16628 31034 16652 31036
rect 16708 31034 16732 31036
rect 16788 31034 16794 31036
rect 16548 30982 16550 31034
rect 16730 30982 16732 31034
rect 16486 30980 16492 30982
rect 16548 30980 16572 30982
rect 16628 30980 16652 30982
rect 16708 30980 16732 30982
rect 16788 30980 16794 30982
rect 16486 30971 16794 30980
rect 9827 30492 10135 30501
rect 9827 30490 9833 30492
rect 9889 30490 9913 30492
rect 9969 30490 9993 30492
rect 10049 30490 10073 30492
rect 10129 30490 10135 30492
rect 9889 30438 9891 30490
rect 10071 30438 10073 30490
rect 9827 30436 9833 30438
rect 9889 30436 9913 30438
rect 9969 30436 9993 30438
rect 10049 30436 10073 30438
rect 10129 30436 10135 30438
rect 9827 30427 10135 30436
rect 14266 30492 14574 30501
rect 14266 30490 14272 30492
rect 14328 30490 14352 30492
rect 14408 30490 14432 30492
rect 14488 30490 14512 30492
rect 14568 30490 14574 30492
rect 14328 30438 14330 30490
rect 14510 30438 14512 30490
rect 14266 30436 14272 30438
rect 14328 30436 14352 30438
rect 14408 30436 14432 30438
rect 14488 30436 14512 30438
rect 14568 30436 14574 30438
rect 14266 30427 14574 30436
rect 18705 30492 19013 30501
rect 18705 30490 18711 30492
rect 18767 30490 18791 30492
rect 18847 30490 18871 30492
rect 18927 30490 18951 30492
rect 19007 30490 19013 30492
rect 18767 30438 18769 30490
rect 18949 30438 18951 30490
rect 18705 30436 18711 30438
rect 18767 30436 18791 30438
rect 18847 30436 18871 30438
rect 18927 30436 18951 30438
rect 19007 30436 19013 30438
rect 18705 30427 19013 30436
rect 8944 30388 8996 30394
rect 8944 30330 8996 30336
rect 8956 28082 8984 30330
rect 12047 29948 12355 29957
rect 12047 29946 12053 29948
rect 12109 29946 12133 29948
rect 12189 29946 12213 29948
rect 12269 29946 12293 29948
rect 12349 29946 12355 29948
rect 12109 29894 12111 29946
rect 12291 29894 12293 29946
rect 12047 29892 12053 29894
rect 12109 29892 12133 29894
rect 12189 29892 12213 29894
rect 12269 29892 12293 29894
rect 12349 29892 12355 29894
rect 12047 29883 12355 29892
rect 16486 29948 16794 29957
rect 16486 29946 16492 29948
rect 16548 29946 16572 29948
rect 16628 29946 16652 29948
rect 16708 29946 16732 29948
rect 16788 29946 16794 29948
rect 16548 29894 16550 29946
rect 16730 29894 16732 29946
rect 16486 29892 16492 29894
rect 16548 29892 16572 29894
rect 16628 29892 16652 29894
rect 16708 29892 16732 29894
rect 16788 29892 16794 29894
rect 16486 29883 16794 29892
rect 9827 29404 10135 29413
rect 9827 29402 9833 29404
rect 9889 29402 9913 29404
rect 9969 29402 9993 29404
rect 10049 29402 10073 29404
rect 10129 29402 10135 29404
rect 9889 29350 9891 29402
rect 10071 29350 10073 29402
rect 9827 29348 9833 29350
rect 9889 29348 9913 29350
rect 9969 29348 9993 29350
rect 10049 29348 10073 29350
rect 10129 29348 10135 29350
rect 9827 29339 10135 29348
rect 14266 29404 14574 29413
rect 14266 29402 14272 29404
rect 14328 29402 14352 29404
rect 14408 29402 14432 29404
rect 14488 29402 14512 29404
rect 14568 29402 14574 29404
rect 14328 29350 14330 29402
rect 14510 29350 14512 29402
rect 14266 29348 14272 29350
rect 14328 29348 14352 29350
rect 14408 29348 14432 29350
rect 14488 29348 14512 29350
rect 14568 29348 14574 29350
rect 14266 29339 14574 29348
rect 18705 29404 19013 29413
rect 18705 29402 18711 29404
rect 18767 29402 18791 29404
rect 18847 29402 18871 29404
rect 18927 29402 18951 29404
rect 19007 29402 19013 29404
rect 18767 29350 18769 29402
rect 18949 29350 18951 29402
rect 18705 29348 18711 29350
rect 18767 29348 18791 29350
rect 18847 29348 18871 29350
rect 18927 29348 18951 29350
rect 19007 29348 19013 29350
rect 18705 29339 19013 29348
rect 12047 28860 12355 28869
rect 12047 28858 12053 28860
rect 12109 28858 12133 28860
rect 12189 28858 12213 28860
rect 12269 28858 12293 28860
rect 12349 28858 12355 28860
rect 12109 28806 12111 28858
rect 12291 28806 12293 28858
rect 12047 28804 12053 28806
rect 12109 28804 12133 28806
rect 12189 28804 12213 28806
rect 12269 28804 12293 28806
rect 12349 28804 12355 28806
rect 12047 28795 12355 28804
rect 16486 28860 16794 28869
rect 16486 28858 16492 28860
rect 16548 28858 16572 28860
rect 16628 28858 16652 28860
rect 16708 28858 16732 28860
rect 16788 28858 16794 28860
rect 16548 28806 16550 28858
rect 16730 28806 16732 28858
rect 16486 28804 16492 28806
rect 16548 28804 16572 28806
rect 16628 28804 16652 28806
rect 16708 28804 16732 28806
rect 16788 28804 16794 28806
rect 16486 28795 16794 28804
rect 9827 28316 10135 28325
rect 9827 28314 9833 28316
rect 9889 28314 9913 28316
rect 9969 28314 9993 28316
rect 10049 28314 10073 28316
rect 10129 28314 10135 28316
rect 9889 28262 9891 28314
rect 10071 28262 10073 28314
rect 9827 28260 9833 28262
rect 9889 28260 9913 28262
rect 9969 28260 9993 28262
rect 10049 28260 10073 28262
rect 10129 28260 10135 28262
rect 9827 28251 10135 28260
rect 14266 28316 14574 28325
rect 14266 28314 14272 28316
rect 14328 28314 14352 28316
rect 14408 28314 14432 28316
rect 14488 28314 14512 28316
rect 14568 28314 14574 28316
rect 14328 28262 14330 28314
rect 14510 28262 14512 28314
rect 14266 28260 14272 28262
rect 14328 28260 14352 28262
rect 14408 28260 14432 28262
rect 14488 28260 14512 28262
rect 14568 28260 14574 28262
rect 14266 28251 14574 28260
rect 18705 28316 19013 28325
rect 18705 28314 18711 28316
rect 18767 28314 18791 28316
rect 18847 28314 18871 28316
rect 18927 28314 18951 28316
rect 19007 28314 19013 28316
rect 18767 28262 18769 28314
rect 18949 28262 18951 28314
rect 18705 28260 18711 28262
rect 18767 28260 18791 28262
rect 18847 28260 18871 28262
rect 18927 28260 18951 28262
rect 19007 28260 19013 28262
rect 18705 28251 19013 28260
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8956 22642 8984 28018
rect 12047 27772 12355 27781
rect 12047 27770 12053 27772
rect 12109 27770 12133 27772
rect 12189 27770 12213 27772
rect 12269 27770 12293 27772
rect 12349 27770 12355 27772
rect 12109 27718 12111 27770
rect 12291 27718 12293 27770
rect 12047 27716 12053 27718
rect 12109 27716 12133 27718
rect 12189 27716 12213 27718
rect 12269 27716 12293 27718
rect 12349 27716 12355 27718
rect 12047 27707 12355 27716
rect 16486 27772 16794 27781
rect 16486 27770 16492 27772
rect 16548 27770 16572 27772
rect 16628 27770 16652 27772
rect 16708 27770 16732 27772
rect 16788 27770 16794 27772
rect 16548 27718 16550 27770
rect 16730 27718 16732 27770
rect 16486 27716 16492 27718
rect 16548 27716 16572 27718
rect 16628 27716 16652 27718
rect 16708 27716 16732 27718
rect 16788 27716 16794 27718
rect 16486 27707 16794 27716
rect 9827 27228 10135 27237
rect 9827 27226 9833 27228
rect 9889 27226 9913 27228
rect 9969 27226 9993 27228
rect 10049 27226 10073 27228
rect 10129 27226 10135 27228
rect 9889 27174 9891 27226
rect 10071 27174 10073 27226
rect 9827 27172 9833 27174
rect 9889 27172 9913 27174
rect 9969 27172 9993 27174
rect 10049 27172 10073 27174
rect 10129 27172 10135 27174
rect 9827 27163 10135 27172
rect 14266 27228 14574 27237
rect 14266 27226 14272 27228
rect 14328 27226 14352 27228
rect 14408 27226 14432 27228
rect 14488 27226 14512 27228
rect 14568 27226 14574 27228
rect 14328 27174 14330 27226
rect 14510 27174 14512 27226
rect 14266 27172 14272 27174
rect 14328 27172 14352 27174
rect 14408 27172 14432 27174
rect 14488 27172 14512 27174
rect 14568 27172 14574 27174
rect 14266 27163 14574 27172
rect 18705 27228 19013 27237
rect 18705 27226 18711 27228
rect 18767 27226 18791 27228
rect 18847 27226 18871 27228
rect 18927 27226 18951 27228
rect 19007 27226 19013 27228
rect 18767 27174 18769 27226
rect 18949 27174 18951 27226
rect 18705 27172 18711 27174
rect 18767 27172 18791 27174
rect 18847 27172 18871 27174
rect 18927 27172 18951 27174
rect 19007 27172 19013 27174
rect 18705 27163 19013 27172
rect 12047 26684 12355 26693
rect 12047 26682 12053 26684
rect 12109 26682 12133 26684
rect 12189 26682 12213 26684
rect 12269 26682 12293 26684
rect 12349 26682 12355 26684
rect 12109 26630 12111 26682
rect 12291 26630 12293 26682
rect 12047 26628 12053 26630
rect 12109 26628 12133 26630
rect 12189 26628 12213 26630
rect 12269 26628 12293 26630
rect 12349 26628 12355 26630
rect 12047 26619 12355 26628
rect 16486 26684 16794 26693
rect 16486 26682 16492 26684
rect 16548 26682 16572 26684
rect 16628 26682 16652 26684
rect 16708 26682 16732 26684
rect 16788 26682 16794 26684
rect 16548 26630 16550 26682
rect 16730 26630 16732 26682
rect 16486 26628 16492 26630
rect 16548 26628 16572 26630
rect 16628 26628 16652 26630
rect 16708 26628 16732 26630
rect 16788 26628 16794 26630
rect 16486 26619 16794 26628
rect 9827 26140 10135 26149
rect 9827 26138 9833 26140
rect 9889 26138 9913 26140
rect 9969 26138 9993 26140
rect 10049 26138 10073 26140
rect 10129 26138 10135 26140
rect 9889 26086 9891 26138
rect 10071 26086 10073 26138
rect 9827 26084 9833 26086
rect 9889 26084 9913 26086
rect 9969 26084 9993 26086
rect 10049 26084 10073 26086
rect 10129 26084 10135 26086
rect 9827 26075 10135 26084
rect 14266 26140 14574 26149
rect 14266 26138 14272 26140
rect 14328 26138 14352 26140
rect 14408 26138 14432 26140
rect 14488 26138 14512 26140
rect 14568 26138 14574 26140
rect 14328 26086 14330 26138
rect 14510 26086 14512 26138
rect 14266 26084 14272 26086
rect 14328 26084 14352 26086
rect 14408 26084 14432 26086
rect 14488 26084 14512 26086
rect 14568 26084 14574 26086
rect 14266 26075 14574 26084
rect 18705 26140 19013 26149
rect 18705 26138 18711 26140
rect 18767 26138 18791 26140
rect 18847 26138 18871 26140
rect 18927 26138 18951 26140
rect 19007 26138 19013 26140
rect 18767 26086 18769 26138
rect 18949 26086 18951 26138
rect 18705 26084 18711 26086
rect 18767 26084 18791 26086
rect 18847 26084 18871 26086
rect 18927 26084 18951 26086
rect 19007 26084 19013 26086
rect 18705 26075 19013 26084
rect 12047 25596 12355 25605
rect 12047 25594 12053 25596
rect 12109 25594 12133 25596
rect 12189 25594 12213 25596
rect 12269 25594 12293 25596
rect 12349 25594 12355 25596
rect 12109 25542 12111 25594
rect 12291 25542 12293 25594
rect 12047 25540 12053 25542
rect 12109 25540 12133 25542
rect 12189 25540 12213 25542
rect 12269 25540 12293 25542
rect 12349 25540 12355 25542
rect 12047 25531 12355 25540
rect 16486 25596 16794 25605
rect 16486 25594 16492 25596
rect 16548 25594 16572 25596
rect 16628 25594 16652 25596
rect 16708 25594 16732 25596
rect 16788 25594 16794 25596
rect 16548 25542 16550 25594
rect 16730 25542 16732 25594
rect 16486 25540 16492 25542
rect 16548 25540 16572 25542
rect 16628 25540 16652 25542
rect 16708 25540 16732 25542
rect 16788 25540 16794 25542
rect 16486 25531 16794 25540
rect 9827 25052 10135 25061
rect 9827 25050 9833 25052
rect 9889 25050 9913 25052
rect 9969 25050 9993 25052
rect 10049 25050 10073 25052
rect 10129 25050 10135 25052
rect 9889 24998 9891 25050
rect 10071 24998 10073 25050
rect 9827 24996 9833 24998
rect 9889 24996 9913 24998
rect 9969 24996 9993 24998
rect 10049 24996 10073 24998
rect 10129 24996 10135 24998
rect 9827 24987 10135 24996
rect 14266 25052 14574 25061
rect 14266 25050 14272 25052
rect 14328 25050 14352 25052
rect 14408 25050 14432 25052
rect 14488 25050 14512 25052
rect 14568 25050 14574 25052
rect 14328 24998 14330 25050
rect 14510 24998 14512 25050
rect 14266 24996 14272 24998
rect 14328 24996 14352 24998
rect 14408 24996 14432 24998
rect 14488 24996 14512 24998
rect 14568 24996 14574 24998
rect 14266 24987 14574 24996
rect 18705 25052 19013 25061
rect 18705 25050 18711 25052
rect 18767 25050 18791 25052
rect 18847 25050 18871 25052
rect 18927 25050 18951 25052
rect 19007 25050 19013 25052
rect 18767 24998 18769 25050
rect 18949 24998 18951 25050
rect 18705 24996 18711 24998
rect 18767 24996 18791 24998
rect 18847 24996 18871 24998
rect 18927 24996 18951 24998
rect 19007 24996 19013 24998
rect 18705 24987 19013 24996
rect 9128 24880 9180 24886
rect 9128 24822 9180 24828
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 8956 21486 8984 22578
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 5388 3227 5696 3236
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 8956 2514 8984 21422
rect 9048 10674 9076 24006
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9140 3738 9168 24822
rect 12047 24508 12355 24517
rect 12047 24506 12053 24508
rect 12109 24506 12133 24508
rect 12189 24506 12213 24508
rect 12269 24506 12293 24508
rect 12349 24506 12355 24508
rect 12109 24454 12111 24506
rect 12291 24454 12293 24506
rect 12047 24452 12053 24454
rect 12109 24452 12133 24454
rect 12189 24452 12213 24454
rect 12269 24452 12293 24454
rect 12349 24452 12355 24454
rect 12047 24443 12355 24452
rect 16486 24508 16794 24517
rect 16486 24506 16492 24508
rect 16548 24506 16572 24508
rect 16628 24506 16652 24508
rect 16708 24506 16732 24508
rect 16788 24506 16794 24508
rect 16548 24454 16550 24506
rect 16730 24454 16732 24506
rect 16486 24452 16492 24454
rect 16548 24452 16572 24454
rect 16628 24452 16652 24454
rect 16708 24452 16732 24454
rect 16788 24452 16794 24454
rect 16486 24443 16794 24452
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9692 6322 9720 24074
rect 9827 23964 10135 23973
rect 9827 23962 9833 23964
rect 9889 23962 9913 23964
rect 9969 23962 9993 23964
rect 10049 23962 10073 23964
rect 10129 23962 10135 23964
rect 9889 23910 9891 23962
rect 10071 23910 10073 23962
rect 9827 23908 9833 23910
rect 9889 23908 9913 23910
rect 9969 23908 9993 23910
rect 10049 23908 10073 23910
rect 10129 23908 10135 23910
rect 9827 23899 10135 23908
rect 14266 23964 14574 23973
rect 14266 23962 14272 23964
rect 14328 23962 14352 23964
rect 14408 23962 14432 23964
rect 14488 23962 14512 23964
rect 14568 23962 14574 23964
rect 14328 23910 14330 23962
rect 14510 23910 14512 23962
rect 14266 23908 14272 23910
rect 14328 23908 14352 23910
rect 14408 23908 14432 23910
rect 14488 23908 14512 23910
rect 14568 23908 14574 23910
rect 14266 23899 14574 23908
rect 18705 23964 19013 23973
rect 18705 23962 18711 23964
rect 18767 23962 18791 23964
rect 18847 23962 18871 23964
rect 18927 23962 18951 23964
rect 19007 23962 19013 23964
rect 18767 23910 18769 23962
rect 18949 23910 18951 23962
rect 18705 23908 18711 23910
rect 18767 23908 18791 23910
rect 18847 23908 18871 23910
rect 18927 23908 18951 23910
rect 19007 23908 19013 23910
rect 18705 23899 19013 23908
rect 12047 23420 12355 23429
rect 12047 23418 12053 23420
rect 12109 23418 12133 23420
rect 12189 23418 12213 23420
rect 12269 23418 12293 23420
rect 12349 23418 12355 23420
rect 12109 23366 12111 23418
rect 12291 23366 12293 23418
rect 12047 23364 12053 23366
rect 12109 23364 12133 23366
rect 12189 23364 12213 23366
rect 12269 23364 12293 23366
rect 12349 23364 12355 23366
rect 12047 23355 12355 23364
rect 16486 23420 16794 23429
rect 16486 23418 16492 23420
rect 16548 23418 16572 23420
rect 16628 23418 16652 23420
rect 16708 23418 16732 23420
rect 16788 23418 16794 23420
rect 16548 23366 16550 23418
rect 16730 23366 16732 23418
rect 16486 23364 16492 23366
rect 16548 23364 16572 23366
rect 16628 23364 16652 23366
rect 16708 23364 16732 23366
rect 16788 23364 16794 23366
rect 16486 23355 16794 23364
rect 9827 22876 10135 22885
rect 9827 22874 9833 22876
rect 9889 22874 9913 22876
rect 9969 22874 9993 22876
rect 10049 22874 10073 22876
rect 10129 22874 10135 22876
rect 9889 22822 9891 22874
rect 10071 22822 10073 22874
rect 9827 22820 9833 22822
rect 9889 22820 9913 22822
rect 9969 22820 9993 22822
rect 10049 22820 10073 22822
rect 10129 22820 10135 22822
rect 9827 22811 10135 22820
rect 14266 22876 14574 22885
rect 14266 22874 14272 22876
rect 14328 22874 14352 22876
rect 14408 22874 14432 22876
rect 14488 22874 14512 22876
rect 14568 22874 14574 22876
rect 14328 22822 14330 22874
rect 14510 22822 14512 22874
rect 14266 22820 14272 22822
rect 14328 22820 14352 22822
rect 14408 22820 14432 22822
rect 14488 22820 14512 22822
rect 14568 22820 14574 22822
rect 14266 22811 14574 22820
rect 18705 22876 19013 22885
rect 18705 22874 18711 22876
rect 18767 22874 18791 22876
rect 18847 22874 18871 22876
rect 18927 22874 18951 22876
rect 19007 22874 19013 22876
rect 18767 22822 18769 22874
rect 18949 22822 18951 22874
rect 18705 22820 18711 22822
rect 18767 22820 18791 22822
rect 18847 22820 18871 22822
rect 18927 22820 18951 22822
rect 19007 22820 19013 22822
rect 18705 22811 19013 22820
rect 12047 22332 12355 22341
rect 12047 22330 12053 22332
rect 12109 22330 12133 22332
rect 12189 22330 12213 22332
rect 12269 22330 12293 22332
rect 12349 22330 12355 22332
rect 12109 22278 12111 22330
rect 12291 22278 12293 22330
rect 12047 22276 12053 22278
rect 12109 22276 12133 22278
rect 12189 22276 12213 22278
rect 12269 22276 12293 22278
rect 12349 22276 12355 22278
rect 12047 22267 12355 22276
rect 16486 22332 16794 22341
rect 16486 22330 16492 22332
rect 16548 22330 16572 22332
rect 16628 22330 16652 22332
rect 16708 22330 16732 22332
rect 16788 22330 16794 22332
rect 16548 22278 16550 22330
rect 16730 22278 16732 22330
rect 16486 22276 16492 22278
rect 16548 22276 16572 22278
rect 16628 22276 16652 22278
rect 16708 22276 16732 22278
rect 16788 22276 16794 22278
rect 16486 22267 16794 22276
rect 9827 21788 10135 21797
rect 9827 21786 9833 21788
rect 9889 21786 9913 21788
rect 9969 21786 9993 21788
rect 10049 21786 10073 21788
rect 10129 21786 10135 21788
rect 9889 21734 9891 21786
rect 10071 21734 10073 21786
rect 9827 21732 9833 21734
rect 9889 21732 9913 21734
rect 9969 21732 9993 21734
rect 10049 21732 10073 21734
rect 10129 21732 10135 21734
rect 9827 21723 10135 21732
rect 14266 21788 14574 21797
rect 14266 21786 14272 21788
rect 14328 21786 14352 21788
rect 14408 21786 14432 21788
rect 14488 21786 14512 21788
rect 14568 21786 14574 21788
rect 14328 21734 14330 21786
rect 14510 21734 14512 21786
rect 14266 21732 14272 21734
rect 14328 21732 14352 21734
rect 14408 21732 14432 21734
rect 14488 21732 14512 21734
rect 14568 21732 14574 21734
rect 14266 21723 14574 21732
rect 18705 21788 19013 21797
rect 18705 21786 18711 21788
rect 18767 21786 18791 21788
rect 18847 21786 18871 21788
rect 18927 21786 18951 21788
rect 19007 21786 19013 21788
rect 18767 21734 18769 21786
rect 18949 21734 18951 21786
rect 18705 21732 18711 21734
rect 18767 21732 18791 21734
rect 18847 21732 18871 21734
rect 18927 21732 18951 21734
rect 19007 21732 19013 21734
rect 18705 21723 19013 21732
rect 12047 21244 12355 21253
rect 12047 21242 12053 21244
rect 12109 21242 12133 21244
rect 12189 21242 12213 21244
rect 12269 21242 12293 21244
rect 12349 21242 12355 21244
rect 12109 21190 12111 21242
rect 12291 21190 12293 21242
rect 12047 21188 12053 21190
rect 12109 21188 12133 21190
rect 12189 21188 12213 21190
rect 12269 21188 12293 21190
rect 12349 21188 12355 21190
rect 12047 21179 12355 21188
rect 16486 21244 16794 21253
rect 16486 21242 16492 21244
rect 16548 21242 16572 21244
rect 16628 21242 16652 21244
rect 16708 21242 16732 21244
rect 16788 21242 16794 21244
rect 16548 21190 16550 21242
rect 16730 21190 16732 21242
rect 16486 21188 16492 21190
rect 16548 21188 16572 21190
rect 16628 21188 16652 21190
rect 16708 21188 16732 21190
rect 16788 21188 16794 21190
rect 16486 21179 16794 21188
rect 9827 20700 10135 20709
rect 9827 20698 9833 20700
rect 9889 20698 9913 20700
rect 9969 20698 9993 20700
rect 10049 20698 10073 20700
rect 10129 20698 10135 20700
rect 9889 20646 9891 20698
rect 10071 20646 10073 20698
rect 9827 20644 9833 20646
rect 9889 20644 9913 20646
rect 9969 20644 9993 20646
rect 10049 20644 10073 20646
rect 10129 20644 10135 20646
rect 9827 20635 10135 20644
rect 14266 20700 14574 20709
rect 14266 20698 14272 20700
rect 14328 20698 14352 20700
rect 14408 20698 14432 20700
rect 14488 20698 14512 20700
rect 14568 20698 14574 20700
rect 14328 20646 14330 20698
rect 14510 20646 14512 20698
rect 14266 20644 14272 20646
rect 14328 20644 14352 20646
rect 14408 20644 14432 20646
rect 14488 20644 14512 20646
rect 14568 20644 14574 20646
rect 14266 20635 14574 20644
rect 18705 20700 19013 20709
rect 18705 20698 18711 20700
rect 18767 20698 18791 20700
rect 18847 20698 18871 20700
rect 18927 20698 18951 20700
rect 19007 20698 19013 20700
rect 18767 20646 18769 20698
rect 18949 20646 18951 20698
rect 18705 20644 18711 20646
rect 18767 20644 18791 20646
rect 18847 20644 18871 20646
rect 18927 20644 18951 20646
rect 19007 20644 19013 20646
rect 18705 20635 19013 20644
rect 12047 20156 12355 20165
rect 12047 20154 12053 20156
rect 12109 20154 12133 20156
rect 12189 20154 12213 20156
rect 12269 20154 12293 20156
rect 12349 20154 12355 20156
rect 12109 20102 12111 20154
rect 12291 20102 12293 20154
rect 12047 20100 12053 20102
rect 12109 20100 12133 20102
rect 12189 20100 12213 20102
rect 12269 20100 12293 20102
rect 12349 20100 12355 20102
rect 12047 20091 12355 20100
rect 16486 20156 16794 20165
rect 16486 20154 16492 20156
rect 16548 20154 16572 20156
rect 16628 20154 16652 20156
rect 16708 20154 16732 20156
rect 16788 20154 16794 20156
rect 16548 20102 16550 20154
rect 16730 20102 16732 20154
rect 16486 20100 16492 20102
rect 16548 20100 16572 20102
rect 16628 20100 16652 20102
rect 16708 20100 16732 20102
rect 16788 20100 16794 20102
rect 16486 20091 16794 20100
rect 9827 19612 10135 19621
rect 9827 19610 9833 19612
rect 9889 19610 9913 19612
rect 9969 19610 9993 19612
rect 10049 19610 10073 19612
rect 10129 19610 10135 19612
rect 9889 19558 9891 19610
rect 10071 19558 10073 19610
rect 9827 19556 9833 19558
rect 9889 19556 9913 19558
rect 9969 19556 9993 19558
rect 10049 19556 10073 19558
rect 10129 19556 10135 19558
rect 9827 19547 10135 19556
rect 14266 19612 14574 19621
rect 14266 19610 14272 19612
rect 14328 19610 14352 19612
rect 14408 19610 14432 19612
rect 14488 19610 14512 19612
rect 14568 19610 14574 19612
rect 14328 19558 14330 19610
rect 14510 19558 14512 19610
rect 14266 19556 14272 19558
rect 14328 19556 14352 19558
rect 14408 19556 14432 19558
rect 14488 19556 14512 19558
rect 14568 19556 14574 19558
rect 14266 19547 14574 19556
rect 18705 19612 19013 19621
rect 18705 19610 18711 19612
rect 18767 19610 18791 19612
rect 18847 19610 18871 19612
rect 18927 19610 18951 19612
rect 19007 19610 19013 19612
rect 18767 19558 18769 19610
rect 18949 19558 18951 19610
rect 18705 19556 18711 19558
rect 18767 19556 18791 19558
rect 18847 19556 18871 19558
rect 18927 19556 18951 19558
rect 19007 19556 19013 19558
rect 18705 19547 19013 19556
rect 12047 19068 12355 19077
rect 12047 19066 12053 19068
rect 12109 19066 12133 19068
rect 12189 19066 12213 19068
rect 12269 19066 12293 19068
rect 12349 19066 12355 19068
rect 12109 19014 12111 19066
rect 12291 19014 12293 19066
rect 12047 19012 12053 19014
rect 12109 19012 12133 19014
rect 12189 19012 12213 19014
rect 12269 19012 12293 19014
rect 12349 19012 12355 19014
rect 12047 19003 12355 19012
rect 16486 19068 16794 19077
rect 16486 19066 16492 19068
rect 16548 19066 16572 19068
rect 16628 19066 16652 19068
rect 16708 19066 16732 19068
rect 16788 19066 16794 19068
rect 16548 19014 16550 19066
rect 16730 19014 16732 19066
rect 16486 19012 16492 19014
rect 16548 19012 16572 19014
rect 16628 19012 16652 19014
rect 16708 19012 16732 19014
rect 16788 19012 16794 19014
rect 16486 19003 16794 19012
rect 9827 18524 10135 18533
rect 9827 18522 9833 18524
rect 9889 18522 9913 18524
rect 9969 18522 9993 18524
rect 10049 18522 10073 18524
rect 10129 18522 10135 18524
rect 9889 18470 9891 18522
rect 10071 18470 10073 18522
rect 9827 18468 9833 18470
rect 9889 18468 9913 18470
rect 9969 18468 9993 18470
rect 10049 18468 10073 18470
rect 10129 18468 10135 18470
rect 9827 18459 10135 18468
rect 14266 18524 14574 18533
rect 14266 18522 14272 18524
rect 14328 18522 14352 18524
rect 14408 18522 14432 18524
rect 14488 18522 14512 18524
rect 14568 18522 14574 18524
rect 14328 18470 14330 18522
rect 14510 18470 14512 18522
rect 14266 18468 14272 18470
rect 14328 18468 14352 18470
rect 14408 18468 14432 18470
rect 14488 18468 14512 18470
rect 14568 18468 14574 18470
rect 14266 18459 14574 18468
rect 18705 18524 19013 18533
rect 18705 18522 18711 18524
rect 18767 18522 18791 18524
rect 18847 18522 18871 18524
rect 18927 18522 18951 18524
rect 19007 18522 19013 18524
rect 18767 18470 18769 18522
rect 18949 18470 18951 18522
rect 18705 18468 18711 18470
rect 18767 18468 18791 18470
rect 18847 18468 18871 18470
rect 18927 18468 18951 18470
rect 19007 18468 19013 18470
rect 18705 18459 19013 18468
rect 12047 17980 12355 17989
rect 12047 17978 12053 17980
rect 12109 17978 12133 17980
rect 12189 17978 12213 17980
rect 12269 17978 12293 17980
rect 12349 17978 12355 17980
rect 12109 17926 12111 17978
rect 12291 17926 12293 17978
rect 12047 17924 12053 17926
rect 12109 17924 12133 17926
rect 12189 17924 12213 17926
rect 12269 17924 12293 17926
rect 12349 17924 12355 17926
rect 12047 17915 12355 17924
rect 16486 17980 16794 17989
rect 16486 17978 16492 17980
rect 16548 17978 16572 17980
rect 16628 17978 16652 17980
rect 16708 17978 16732 17980
rect 16788 17978 16794 17980
rect 16548 17926 16550 17978
rect 16730 17926 16732 17978
rect 16486 17924 16492 17926
rect 16548 17924 16572 17926
rect 16628 17924 16652 17926
rect 16708 17924 16732 17926
rect 16788 17924 16794 17926
rect 16486 17915 16794 17924
rect 9827 17436 10135 17445
rect 9827 17434 9833 17436
rect 9889 17434 9913 17436
rect 9969 17434 9993 17436
rect 10049 17434 10073 17436
rect 10129 17434 10135 17436
rect 9889 17382 9891 17434
rect 10071 17382 10073 17434
rect 9827 17380 9833 17382
rect 9889 17380 9913 17382
rect 9969 17380 9993 17382
rect 10049 17380 10073 17382
rect 10129 17380 10135 17382
rect 9827 17371 10135 17380
rect 14266 17436 14574 17445
rect 14266 17434 14272 17436
rect 14328 17434 14352 17436
rect 14408 17434 14432 17436
rect 14488 17434 14512 17436
rect 14568 17434 14574 17436
rect 14328 17382 14330 17434
rect 14510 17382 14512 17434
rect 14266 17380 14272 17382
rect 14328 17380 14352 17382
rect 14408 17380 14432 17382
rect 14488 17380 14512 17382
rect 14568 17380 14574 17382
rect 14266 17371 14574 17380
rect 18705 17436 19013 17445
rect 18705 17434 18711 17436
rect 18767 17434 18791 17436
rect 18847 17434 18871 17436
rect 18927 17434 18951 17436
rect 19007 17434 19013 17436
rect 18767 17382 18769 17434
rect 18949 17382 18951 17434
rect 18705 17380 18711 17382
rect 18767 17380 18791 17382
rect 18847 17380 18871 17382
rect 18927 17380 18951 17382
rect 19007 17380 19013 17382
rect 18705 17371 19013 17380
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 9827 16348 10135 16357
rect 9827 16346 9833 16348
rect 9889 16346 9913 16348
rect 9969 16346 9993 16348
rect 10049 16346 10073 16348
rect 10129 16346 10135 16348
rect 9889 16294 9891 16346
rect 10071 16294 10073 16346
rect 9827 16292 9833 16294
rect 9889 16292 9913 16294
rect 9969 16292 9993 16294
rect 10049 16292 10073 16294
rect 10129 16292 10135 16294
rect 9827 16283 10135 16292
rect 14266 16348 14574 16357
rect 14266 16346 14272 16348
rect 14328 16346 14352 16348
rect 14408 16346 14432 16348
rect 14488 16346 14512 16348
rect 14568 16346 14574 16348
rect 14328 16294 14330 16346
rect 14510 16294 14512 16346
rect 14266 16292 14272 16294
rect 14328 16292 14352 16294
rect 14408 16292 14432 16294
rect 14488 16292 14512 16294
rect 14568 16292 14574 16294
rect 14266 16283 14574 16292
rect 18705 16348 19013 16357
rect 18705 16346 18711 16348
rect 18767 16346 18791 16348
rect 18847 16346 18871 16348
rect 18927 16346 18951 16348
rect 19007 16346 19013 16348
rect 18767 16294 18769 16346
rect 18949 16294 18951 16346
rect 18705 16292 18711 16294
rect 18767 16292 18791 16294
rect 18847 16292 18871 16294
rect 18927 16292 18951 16294
rect 19007 16292 19013 16294
rect 18705 16283 19013 16292
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 9827 15260 10135 15269
rect 9827 15258 9833 15260
rect 9889 15258 9913 15260
rect 9969 15258 9993 15260
rect 10049 15258 10073 15260
rect 10129 15258 10135 15260
rect 9889 15206 9891 15258
rect 10071 15206 10073 15258
rect 9827 15204 9833 15206
rect 9889 15204 9913 15206
rect 9969 15204 9993 15206
rect 10049 15204 10073 15206
rect 10129 15204 10135 15206
rect 9827 15195 10135 15204
rect 14266 15260 14574 15269
rect 14266 15258 14272 15260
rect 14328 15258 14352 15260
rect 14408 15258 14432 15260
rect 14488 15258 14512 15260
rect 14568 15258 14574 15260
rect 14328 15206 14330 15258
rect 14510 15206 14512 15258
rect 14266 15204 14272 15206
rect 14328 15204 14352 15206
rect 14408 15204 14432 15206
rect 14488 15204 14512 15206
rect 14568 15204 14574 15206
rect 14266 15195 14574 15204
rect 18705 15260 19013 15269
rect 18705 15258 18711 15260
rect 18767 15258 18791 15260
rect 18847 15258 18871 15260
rect 18927 15258 18951 15260
rect 19007 15258 19013 15260
rect 18767 15206 18769 15258
rect 18949 15206 18951 15258
rect 18705 15204 18711 15206
rect 18767 15204 18791 15206
rect 18847 15204 18871 15206
rect 18927 15204 18951 15206
rect 19007 15204 19013 15206
rect 18705 15195 19013 15204
rect 12047 14716 12355 14725
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 9827 14172 10135 14181
rect 9827 14170 9833 14172
rect 9889 14170 9913 14172
rect 9969 14170 9993 14172
rect 10049 14170 10073 14172
rect 10129 14170 10135 14172
rect 9889 14118 9891 14170
rect 10071 14118 10073 14170
rect 9827 14116 9833 14118
rect 9889 14116 9913 14118
rect 9969 14116 9993 14118
rect 10049 14116 10073 14118
rect 10129 14116 10135 14118
rect 9827 14107 10135 14116
rect 14266 14172 14574 14181
rect 14266 14170 14272 14172
rect 14328 14170 14352 14172
rect 14408 14170 14432 14172
rect 14488 14170 14512 14172
rect 14568 14170 14574 14172
rect 14328 14118 14330 14170
rect 14510 14118 14512 14170
rect 14266 14116 14272 14118
rect 14328 14116 14352 14118
rect 14408 14116 14432 14118
rect 14488 14116 14512 14118
rect 14568 14116 14574 14118
rect 14266 14107 14574 14116
rect 18705 14172 19013 14181
rect 18705 14170 18711 14172
rect 18767 14170 18791 14172
rect 18847 14170 18871 14172
rect 18927 14170 18951 14172
rect 19007 14170 19013 14172
rect 18767 14118 18769 14170
rect 18949 14118 18951 14170
rect 18705 14116 18711 14118
rect 18767 14116 18791 14118
rect 18847 14116 18871 14118
rect 18927 14116 18951 14118
rect 19007 14116 19013 14118
rect 18705 14107 19013 14116
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 9827 13084 10135 13093
rect 9827 13082 9833 13084
rect 9889 13082 9913 13084
rect 9969 13082 9993 13084
rect 10049 13082 10073 13084
rect 10129 13082 10135 13084
rect 9889 13030 9891 13082
rect 10071 13030 10073 13082
rect 9827 13028 9833 13030
rect 9889 13028 9913 13030
rect 9969 13028 9993 13030
rect 10049 13028 10073 13030
rect 10129 13028 10135 13030
rect 9827 13019 10135 13028
rect 14266 13084 14574 13093
rect 14266 13082 14272 13084
rect 14328 13082 14352 13084
rect 14408 13082 14432 13084
rect 14488 13082 14512 13084
rect 14568 13082 14574 13084
rect 14328 13030 14330 13082
rect 14510 13030 14512 13082
rect 14266 13028 14272 13030
rect 14328 13028 14352 13030
rect 14408 13028 14432 13030
rect 14488 13028 14512 13030
rect 14568 13028 14574 13030
rect 14266 13019 14574 13028
rect 18705 13084 19013 13093
rect 18705 13082 18711 13084
rect 18767 13082 18791 13084
rect 18847 13082 18871 13084
rect 18927 13082 18951 13084
rect 19007 13082 19013 13084
rect 18767 13030 18769 13082
rect 18949 13030 18951 13082
rect 18705 13028 18711 13030
rect 18767 13028 18791 13030
rect 18847 13028 18871 13030
rect 18927 13028 18951 13030
rect 19007 13028 19013 13030
rect 18705 13019 19013 13028
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 9827 11996 10135 12005
rect 9827 11994 9833 11996
rect 9889 11994 9913 11996
rect 9969 11994 9993 11996
rect 10049 11994 10073 11996
rect 10129 11994 10135 11996
rect 9889 11942 9891 11994
rect 10071 11942 10073 11994
rect 9827 11940 9833 11942
rect 9889 11940 9913 11942
rect 9969 11940 9993 11942
rect 10049 11940 10073 11942
rect 10129 11940 10135 11942
rect 9827 11931 10135 11940
rect 14266 11996 14574 12005
rect 14266 11994 14272 11996
rect 14328 11994 14352 11996
rect 14408 11994 14432 11996
rect 14488 11994 14512 11996
rect 14568 11994 14574 11996
rect 14328 11942 14330 11994
rect 14510 11942 14512 11994
rect 14266 11940 14272 11942
rect 14328 11940 14352 11942
rect 14408 11940 14432 11942
rect 14488 11940 14512 11942
rect 14568 11940 14574 11942
rect 14266 11931 14574 11940
rect 18705 11996 19013 12005
rect 18705 11994 18711 11996
rect 18767 11994 18791 11996
rect 18847 11994 18871 11996
rect 18927 11994 18951 11996
rect 19007 11994 19013 11996
rect 18767 11942 18769 11994
rect 18949 11942 18951 11994
rect 18705 11940 18711 11942
rect 18767 11940 18791 11942
rect 18847 11940 18871 11942
rect 18927 11940 18951 11942
rect 19007 11940 19013 11942
rect 18705 11931 19013 11940
rect 12047 11452 12355 11461
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 9827 10908 10135 10917
rect 9827 10906 9833 10908
rect 9889 10906 9913 10908
rect 9969 10906 9993 10908
rect 10049 10906 10073 10908
rect 10129 10906 10135 10908
rect 9889 10854 9891 10906
rect 10071 10854 10073 10906
rect 9827 10852 9833 10854
rect 9889 10852 9913 10854
rect 9969 10852 9993 10854
rect 10049 10852 10073 10854
rect 10129 10852 10135 10854
rect 9827 10843 10135 10852
rect 14266 10908 14574 10917
rect 14266 10906 14272 10908
rect 14328 10906 14352 10908
rect 14408 10906 14432 10908
rect 14488 10906 14512 10908
rect 14568 10906 14574 10908
rect 14328 10854 14330 10906
rect 14510 10854 14512 10906
rect 14266 10852 14272 10854
rect 14328 10852 14352 10854
rect 14408 10852 14432 10854
rect 14488 10852 14512 10854
rect 14568 10852 14574 10854
rect 14266 10843 14574 10852
rect 18705 10908 19013 10917
rect 18705 10906 18711 10908
rect 18767 10906 18791 10908
rect 18847 10906 18871 10908
rect 18927 10906 18951 10908
rect 19007 10906 19013 10908
rect 18767 10854 18769 10906
rect 18949 10854 18951 10906
rect 18705 10852 18711 10854
rect 18767 10852 18791 10854
rect 18847 10852 18871 10854
rect 18927 10852 18951 10854
rect 19007 10852 19013 10854
rect 18705 10843 19013 10852
rect 12047 10364 12355 10373
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 16486 10364 16794 10373
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 9827 9820 10135 9829
rect 9827 9818 9833 9820
rect 9889 9818 9913 9820
rect 9969 9818 9993 9820
rect 10049 9818 10073 9820
rect 10129 9818 10135 9820
rect 9889 9766 9891 9818
rect 10071 9766 10073 9818
rect 9827 9764 9833 9766
rect 9889 9764 9913 9766
rect 9969 9764 9993 9766
rect 10049 9764 10073 9766
rect 10129 9764 10135 9766
rect 9827 9755 10135 9764
rect 14266 9820 14574 9829
rect 14266 9818 14272 9820
rect 14328 9818 14352 9820
rect 14408 9818 14432 9820
rect 14488 9818 14512 9820
rect 14568 9818 14574 9820
rect 14328 9766 14330 9818
rect 14510 9766 14512 9818
rect 14266 9764 14272 9766
rect 14328 9764 14352 9766
rect 14408 9764 14432 9766
rect 14488 9764 14512 9766
rect 14568 9764 14574 9766
rect 14266 9755 14574 9764
rect 18705 9820 19013 9829
rect 18705 9818 18711 9820
rect 18767 9818 18791 9820
rect 18847 9818 18871 9820
rect 18927 9818 18951 9820
rect 19007 9818 19013 9820
rect 18767 9766 18769 9818
rect 18949 9766 18951 9818
rect 18705 9764 18711 9766
rect 18767 9764 18791 9766
rect 18847 9764 18871 9766
rect 18927 9764 18951 9766
rect 19007 9764 19013 9766
rect 18705 9755 19013 9764
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 9827 8732 10135 8741
rect 9827 8730 9833 8732
rect 9889 8730 9913 8732
rect 9969 8730 9993 8732
rect 10049 8730 10073 8732
rect 10129 8730 10135 8732
rect 9889 8678 9891 8730
rect 10071 8678 10073 8730
rect 9827 8676 9833 8678
rect 9889 8676 9913 8678
rect 9969 8676 9993 8678
rect 10049 8676 10073 8678
rect 10129 8676 10135 8678
rect 9827 8667 10135 8676
rect 14266 8732 14574 8741
rect 14266 8730 14272 8732
rect 14328 8730 14352 8732
rect 14408 8730 14432 8732
rect 14488 8730 14512 8732
rect 14568 8730 14574 8732
rect 14328 8678 14330 8730
rect 14510 8678 14512 8730
rect 14266 8676 14272 8678
rect 14328 8676 14352 8678
rect 14408 8676 14432 8678
rect 14488 8676 14512 8678
rect 14568 8676 14574 8678
rect 14266 8667 14574 8676
rect 18705 8732 19013 8741
rect 18705 8730 18711 8732
rect 18767 8730 18791 8732
rect 18847 8730 18871 8732
rect 18927 8730 18951 8732
rect 19007 8730 19013 8732
rect 18767 8678 18769 8730
rect 18949 8678 18951 8730
rect 18705 8676 18711 8678
rect 18767 8676 18791 8678
rect 18847 8676 18871 8678
rect 18927 8676 18951 8678
rect 19007 8676 19013 8678
rect 18705 8667 19013 8676
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 14936 800 14964 2382
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 4986 0 5042 800
rect 14922 0 14978 800
<< via2 >>
rect 938 47912 994 47968
rect 3175 47354 3231 47356
rect 3255 47354 3311 47356
rect 3335 47354 3391 47356
rect 3415 47354 3471 47356
rect 3175 47302 3221 47354
rect 3221 47302 3231 47354
rect 3255 47302 3285 47354
rect 3285 47302 3297 47354
rect 3297 47302 3311 47354
rect 3335 47302 3349 47354
rect 3349 47302 3361 47354
rect 3361 47302 3391 47354
rect 3415 47302 3425 47354
rect 3425 47302 3471 47354
rect 3175 47300 3231 47302
rect 3255 47300 3311 47302
rect 3335 47300 3391 47302
rect 3415 47300 3471 47302
rect 7614 47354 7670 47356
rect 7694 47354 7750 47356
rect 7774 47354 7830 47356
rect 7854 47354 7910 47356
rect 7614 47302 7660 47354
rect 7660 47302 7670 47354
rect 7694 47302 7724 47354
rect 7724 47302 7736 47354
rect 7736 47302 7750 47354
rect 7774 47302 7788 47354
rect 7788 47302 7800 47354
rect 7800 47302 7830 47354
rect 7854 47302 7864 47354
rect 7864 47302 7910 47354
rect 7614 47300 7670 47302
rect 7694 47300 7750 47302
rect 7774 47300 7830 47302
rect 7854 47300 7910 47302
rect 12053 47354 12109 47356
rect 12133 47354 12189 47356
rect 12213 47354 12269 47356
rect 12293 47354 12349 47356
rect 12053 47302 12099 47354
rect 12099 47302 12109 47354
rect 12133 47302 12163 47354
rect 12163 47302 12175 47354
rect 12175 47302 12189 47354
rect 12213 47302 12227 47354
rect 12227 47302 12239 47354
rect 12239 47302 12269 47354
rect 12293 47302 12303 47354
rect 12303 47302 12349 47354
rect 12053 47300 12109 47302
rect 12133 47300 12189 47302
rect 12213 47300 12269 47302
rect 12293 47300 12349 47302
rect 16492 47354 16548 47356
rect 16572 47354 16628 47356
rect 16652 47354 16708 47356
rect 16732 47354 16788 47356
rect 16492 47302 16538 47354
rect 16538 47302 16548 47354
rect 16572 47302 16602 47354
rect 16602 47302 16614 47354
rect 16614 47302 16628 47354
rect 16652 47302 16666 47354
rect 16666 47302 16678 47354
rect 16678 47302 16708 47354
rect 16732 47302 16742 47354
rect 16742 47302 16788 47354
rect 16492 47300 16548 47302
rect 16572 47300 16628 47302
rect 16652 47300 16708 47302
rect 16732 47300 16788 47302
rect 938 44376 994 44432
rect 938 40840 994 40896
rect 938 37304 994 37360
rect 938 33768 994 33824
rect 938 30232 994 30288
rect 938 26696 994 26752
rect 938 23160 994 23216
rect 938 19624 994 19680
rect 938 16088 994 16144
rect 938 12552 994 12608
rect 5394 46810 5450 46812
rect 5474 46810 5530 46812
rect 5554 46810 5610 46812
rect 5634 46810 5690 46812
rect 5394 46758 5440 46810
rect 5440 46758 5450 46810
rect 5474 46758 5504 46810
rect 5504 46758 5516 46810
rect 5516 46758 5530 46810
rect 5554 46758 5568 46810
rect 5568 46758 5580 46810
rect 5580 46758 5610 46810
rect 5634 46758 5644 46810
rect 5644 46758 5690 46810
rect 5394 46756 5450 46758
rect 5474 46756 5530 46758
rect 5554 46756 5610 46758
rect 5634 46756 5690 46758
rect 9833 46810 9889 46812
rect 9913 46810 9969 46812
rect 9993 46810 10049 46812
rect 10073 46810 10129 46812
rect 9833 46758 9879 46810
rect 9879 46758 9889 46810
rect 9913 46758 9943 46810
rect 9943 46758 9955 46810
rect 9955 46758 9969 46810
rect 9993 46758 10007 46810
rect 10007 46758 10019 46810
rect 10019 46758 10049 46810
rect 10073 46758 10083 46810
rect 10083 46758 10129 46810
rect 9833 46756 9889 46758
rect 9913 46756 9969 46758
rect 9993 46756 10049 46758
rect 10073 46756 10129 46758
rect 14272 46810 14328 46812
rect 14352 46810 14408 46812
rect 14432 46810 14488 46812
rect 14512 46810 14568 46812
rect 14272 46758 14318 46810
rect 14318 46758 14328 46810
rect 14352 46758 14382 46810
rect 14382 46758 14394 46810
rect 14394 46758 14408 46810
rect 14432 46758 14446 46810
rect 14446 46758 14458 46810
rect 14458 46758 14488 46810
rect 14512 46758 14522 46810
rect 14522 46758 14568 46810
rect 14272 46756 14328 46758
rect 14352 46756 14408 46758
rect 14432 46756 14488 46758
rect 14512 46756 14568 46758
rect 18711 46810 18767 46812
rect 18791 46810 18847 46812
rect 18871 46810 18927 46812
rect 18951 46810 19007 46812
rect 18711 46758 18757 46810
rect 18757 46758 18767 46810
rect 18791 46758 18821 46810
rect 18821 46758 18833 46810
rect 18833 46758 18847 46810
rect 18871 46758 18885 46810
rect 18885 46758 18897 46810
rect 18897 46758 18927 46810
rect 18951 46758 18961 46810
rect 18961 46758 19007 46810
rect 18711 46756 18767 46758
rect 18791 46756 18847 46758
rect 18871 46756 18927 46758
rect 18951 46756 19007 46758
rect 3175 46266 3231 46268
rect 3255 46266 3311 46268
rect 3335 46266 3391 46268
rect 3415 46266 3471 46268
rect 3175 46214 3221 46266
rect 3221 46214 3231 46266
rect 3255 46214 3285 46266
rect 3285 46214 3297 46266
rect 3297 46214 3311 46266
rect 3335 46214 3349 46266
rect 3349 46214 3361 46266
rect 3361 46214 3391 46266
rect 3415 46214 3425 46266
rect 3425 46214 3471 46266
rect 3175 46212 3231 46214
rect 3255 46212 3311 46214
rect 3335 46212 3391 46214
rect 3415 46212 3471 46214
rect 7614 46266 7670 46268
rect 7694 46266 7750 46268
rect 7774 46266 7830 46268
rect 7854 46266 7910 46268
rect 7614 46214 7660 46266
rect 7660 46214 7670 46266
rect 7694 46214 7724 46266
rect 7724 46214 7736 46266
rect 7736 46214 7750 46266
rect 7774 46214 7788 46266
rect 7788 46214 7800 46266
rect 7800 46214 7830 46266
rect 7854 46214 7864 46266
rect 7864 46214 7910 46266
rect 7614 46212 7670 46214
rect 7694 46212 7750 46214
rect 7774 46212 7830 46214
rect 7854 46212 7910 46214
rect 12053 46266 12109 46268
rect 12133 46266 12189 46268
rect 12213 46266 12269 46268
rect 12293 46266 12349 46268
rect 12053 46214 12099 46266
rect 12099 46214 12109 46266
rect 12133 46214 12163 46266
rect 12163 46214 12175 46266
rect 12175 46214 12189 46266
rect 12213 46214 12227 46266
rect 12227 46214 12239 46266
rect 12239 46214 12269 46266
rect 12293 46214 12303 46266
rect 12303 46214 12349 46266
rect 12053 46212 12109 46214
rect 12133 46212 12189 46214
rect 12213 46212 12269 46214
rect 12293 46212 12349 46214
rect 16492 46266 16548 46268
rect 16572 46266 16628 46268
rect 16652 46266 16708 46268
rect 16732 46266 16788 46268
rect 16492 46214 16538 46266
rect 16538 46214 16548 46266
rect 16572 46214 16602 46266
rect 16602 46214 16614 46266
rect 16614 46214 16628 46266
rect 16652 46214 16666 46266
rect 16666 46214 16678 46266
rect 16678 46214 16708 46266
rect 16732 46214 16742 46266
rect 16742 46214 16788 46266
rect 16492 46212 16548 46214
rect 16572 46212 16628 46214
rect 16652 46212 16708 46214
rect 16732 46212 16788 46214
rect 5394 45722 5450 45724
rect 5474 45722 5530 45724
rect 5554 45722 5610 45724
rect 5634 45722 5690 45724
rect 5394 45670 5440 45722
rect 5440 45670 5450 45722
rect 5474 45670 5504 45722
rect 5504 45670 5516 45722
rect 5516 45670 5530 45722
rect 5554 45670 5568 45722
rect 5568 45670 5580 45722
rect 5580 45670 5610 45722
rect 5634 45670 5644 45722
rect 5644 45670 5690 45722
rect 5394 45668 5450 45670
rect 5474 45668 5530 45670
rect 5554 45668 5610 45670
rect 5634 45668 5690 45670
rect 9833 45722 9889 45724
rect 9913 45722 9969 45724
rect 9993 45722 10049 45724
rect 10073 45722 10129 45724
rect 9833 45670 9879 45722
rect 9879 45670 9889 45722
rect 9913 45670 9943 45722
rect 9943 45670 9955 45722
rect 9955 45670 9969 45722
rect 9993 45670 10007 45722
rect 10007 45670 10019 45722
rect 10019 45670 10049 45722
rect 10073 45670 10083 45722
rect 10083 45670 10129 45722
rect 9833 45668 9889 45670
rect 9913 45668 9969 45670
rect 9993 45668 10049 45670
rect 10073 45668 10129 45670
rect 14272 45722 14328 45724
rect 14352 45722 14408 45724
rect 14432 45722 14488 45724
rect 14512 45722 14568 45724
rect 14272 45670 14318 45722
rect 14318 45670 14328 45722
rect 14352 45670 14382 45722
rect 14382 45670 14394 45722
rect 14394 45670 14408 45722
rect 14432 45670 14446 45722
rect 14446 45670 14458 45722
rect 14458 45670 14488 45722
rect 14512 45670 14522 45722
rect 14522 45670 14568 45722
rect 14272 45668 14328 45670
rect 14352 45668 14408 45670
rect 14432 45668 14488 45670
rect 14512 45668 14568 45670
rect 18711 45722 18767 45724
rect 18791 45722 18847 45724
rect 18871 45722 18927 45724
rect 18951 45722 19007 45724
rect 18711 45670 18757 45722
rect 18757 45670 18767 45722
rect 18791 45670 18821 45722
rect 18821 45670 18833 45722
rect 18833 45670 18847 45722
rect 18871 45670 18885 45722
rect 18885 45670 18897 45722
rect 18897 45670 18927 45722
rect 18951 45670 18961 45722
rect 18961 45670 19007 45722
rect 18711 45668 18767 45670
rect 18791 45668 18847 45670
rect 18871 45668 18927 45670
rect 18951 45668 19007 45670
rect 3175 45178 3231 45180
rect 3255 45178 3311 45180
rect 3335 45178 3391 45180
rect 3415 45178 3471 45180
rect 3175 45126 3221 45178
rect 3221 45126 3231 45178
rect 3255 45126 3285 45178
rect 3285 45126 3297 45178
rect 3297 45126 3311 45178
rect 3335 45126 3349 45178
rect 3349 45126 3361 45178
rect 3361 45126 3391 45178
rect 3415 45126 3425 45178
rect 3425 45126 3471 45178
rect 3175 45124 3231 45126
rect 3255 45124 3311 45126
rect 3335 45124 3391 45126
rect 3415 45124 3471 45126
rect 7614 45178 7670 45180
rect 7694 45178 7750 45180
rect 7774 45178 7830 45180
rect 7854 45178 7910 45180
rect 7614 45126 7660 45178
rect 7660 45126 7670 45178
rect 7694 45126 7724 45178
rect 7724 45126 7736 45178
rect 7736 45126 7750 45178
rect 7774 45126 7788 45178
rect 7788 45126 7800 45178
rect 7800 45126 7830 45178
rect 7854 45126 7864 45178
rect 7864 45126 7910 45178
rect 7614 45124 7670 45126
rect 7694 45124 7750 45126
rect 7774 45124 7830 45126
rect 7854 45124 7910 45126
rect 12053 45178 12109 45180
rect 12133 45178 12189 45180
rect 12213 45178 12269 45180
rect 12293 45178 12349 45180
rect 12053 45126 12099 45178
rect 12099 45126 12109 45178
rect 12133 45126 12163 45178
rect 12163 45126 12175 45178
rect 12175 45126 12189 45178
rect 12213 45126 12227 45178
rect 12227 45126 12239 45178
rect 12239 45126 12269 45178
rect 12293 45126 12303 45178
rect 12303 45126 12349 45178
rect 12053 45124 12109 45126
rect 12133 45124 12189 45126
rect 12213 45124 12269 45126
rect 12293 45124 12349 45126
rect 16492 45178 16548 45180
rect 16572 45178 16628 45180
rect 16652 45178 16708 45180
rect 16732 45178 16788 45180
rect 16492 45126 16538 45178
rect 16538 45126 16548 45178
rect 16572 45126 16602 45178
rect 16602 45126 16614 45178
rect 16614 45126 16628 45178
rect 16652 45126 16666 45178
rect 16666 45126 16678 45178
rect 16678 45126 16708 45178
rect 16732 45126 16742 45178
rect 16742 45126 16788 45178
rect 16492 45124 16548 45126
rect 16572 45124 16628 45126
rect 16652 45124 16708 45126
rect 16732 45124 16788 45126
rect 5394 44634 5450 44636
rect 5474 44634 5530 44636
rect 5554 44634 5610 44636
rect 5634 44634 5690 44636
rect 5394 44582 5440 44634
rect 5440 44582 5450 44634
rect 5474 44582 5504 44634
rect 5504 44582 5516 44634
rect 5516 44582 5530 44634
rect 5554 44582 5568 44634
rect 5568 44582 5580 44634
rect 5580 44582 5610 44634
rect 5634 44582 5644 44634
rect 5644 44582 5690 44634
rect 5394 44580 5450 44582
rect 5474 44580 5530 44582
rect 5554 44580 5610 44582
rect 5634 44580 5690 44582
rect 9833 44634 9889 44636
rect 9913 44634 9969 44636
rect 9993 44634 10049 44636
rect 10073 44634 10129 44636
rect 9833 44582 9879 44634
rect 9879 44582 9889 44634
rect 9913 44582 9943 44634
rect 9943 44582 9955 44634
rect 9955 44582 9969 44634
rect 9993 44582 10007 44634
rect 10007 44582 10019 44634
rect 10019 44582 10049 44634
rect 10073 44582 10083 44634
rect 10083 44582 10129 44634
rect 9833 44580 9889 44582
rect 9913 44580 9969 44582
rect 9993 44580 10049 44582
rect 10073 44580 10129 44582
rect 14272 44634 14328 44636
rect 14352 44634 14408 44636
rect 14432 44634 14488 44636
rect 14512 44634 14568 44636
rect 14272 44582 14318 44634
rect 14318 44582 14328 44634
rect 14352 44582 14382 44634
rect 14382 44582 14394 44634
rect 14394 44582 14408 44634
rect 14432 44582 14446 44634
rect 14446 44582 14458 44634
rect 14458 44582 14488 44634
rect 14512 44582 14522 44634
rect 14522 44582 14568 44634
rect 14272 44580 14328 44582
rect 14352 44580 14408 44582
rect 14432 44580 14488 44582
rect 14512 44580 14568 44582
rect 18711 44634 18767 44636
rect 18791 44634 18847 44636
rect 18871 44634 18927 44636
rect 18951 44634 19007 44636
rect 18711 44582 18757 44634
rect 18757 44582 18767 44634
rect 18791 44582 18821 44634
rect 18821 44582 18833 44634
rect 18833 44582 18847 44634
rect 18871 44582 18885 44634
rect 18885 44582 18897 44634
rect 18897 44582 18927 44634
rect 18951 44582 18961 44634
rect 18961 44582 19007 44634
rect 18711 44580 18767 44582
rect 18791 44580 18847 44582
rect 18871 44580 18927 44582
rect 18951 44580 19007 44582
rect 3175 44090 3231 44092
rect 3255 44090 3311 44092
rect 3335 44090 3391 44092
rect 3415 44090 3471 44092
rect 3175 44038 3221 44090
rect 3221 44038 3231 44090
rect 3255 44038 3285 44090
rect 3285 44038 3297 44090
rect 3297 44038 3311 44090
rect 3335 44038 3349 44090
rect 3349 44038 3361 44090
rect 3361 44038 3391 44090
rect 3415 44038 3425 44090
rect 3425 44038 3471 44090
rect 3175 44036 3231 44038
rect 3255 44036 3311 44038
rect 3335 44036 3391 44038
rect 3415 44036 3471 44038
rect 7614 44090 7670 44092
rect 7694 44090 7750 44092
rect 7774 44090 7830 44092
rect 7854 44090 7910 44092
rect 7614 44038 7660 44090
rect 7660 44038 7670 44090
rect 7694 44038 7724 44090
rect 7724 44038 7736 44090
rect 7736 44038 7750 44090
rect 7774 44038 7788 44090
rect 7788 44038 7800 44090
rect 7800 44038 7830 44090
rect 7854 44038 7864 44090
rect 7864 44038 7910 44090
rect 7614 44036 7670 44038
rect 7694 44036 7750 44038
rect 7774 44036 7830 44038
rect 7854 44036 7910 44038
rect 12053 44090 12109 44092
rect 12133 44090 12189 44092
rect 12213 44090 12269 44092
rect 12293 44090 12349 44092
rect 12053 44038 12099 44090
rect 12099 44038 12109 44090
rect 12133 44038 12163 44090
rect 12163 44038 12175 44090
rect 12175 44038 12189 44090
rect 12213 44038 12227 44090
rect 12227 44038 12239 44090
rect 12239 44038 12269 44090
rect 12293 44038 12303 44090
rect 12303 44038 12349 44090
rect 12053 44036 12109 44038
rect 12133 44036 12189 44038
rect 12213 44036 12269 44038
rect 12293 44036 12349 44038
rect 16492 44090 16548 44092
rect 16572 44090 16628 44092
rect 16652 44090 16708 44092
rect 16732 44090 16788 44092
rect 16492 44038 16538 44090
rect 16538 44038 16548 44090
rect 16572 44038 16602 44090
rect 16602 44038 16614 44090
rect 16614 44038 16628 44090
rect 16652 44038 16666 44090
rect 16666 44038 16678 44090
rect 16678 44038 16708 44090
rect 16732 44038 16742 44090
rect 16742 44038 16788 44090
rect 16492 44036 16548 44038
rect 16572 44036 16628 44038
rect 16652 44036 16708 44038
rect 16732 44036 16788 44038
rect 5394 43546 5450 43548
rect 5474 43546 5530 43548
rect 5554 43546 5610 43548
rect 5634 43546 5690 43548
rect 5394 43494 5440 43546
rect 5440 43494 5450 43546
rect 5474 43494 5504 43546
rect 5504 43494 5516 43546
rect 5516 43494 5530 43546
rect 5554 43494 5568 43546
rect 5568 43494 5580 43546
rect 5580 43494 5610 43546
rect 5634 43494 5644 43546
rect 5644 43494 5690 43546
rect 5394 43492 5450 43494
rect 5474 43492 5530 43494
rect 5554 43492 5610 43494
rect 5634 43492 5690 43494
rect 9833 43546 9889 43548
rect 9913 43546 9969 43548
rect 9993 43546 10049 43548
rect 10073 43546 10129 43548
rect 9833 43494 9879 43546
rect 9879 43494 9889 43546
rect 9913 43494 9943 43546
rect 9943 43494 9955 43546
rect 9955 43494 9969 43546
rect 9993 43494 10007 43546
rect 10007 43494 10019 43546
rect 10019 43494 10049 43546
rect 10073 43494 10083 43546
rect 10083 43494 10129 43546
rect 9833 43492 9889 43494
rect 9913 43492 9969 43494
rect 9993 43492 10049 43494
rect 10073 43492 10129 43494
rect 14272 43546 14328 43548
rect 14352 43546 14408 43548
rect 14432 43546 14488 43548
rect 14512 43546 14568 43548
rect 14272 43494 14318 43546
rect 14318 43494 14328 43546
rect 14352 43494 14382 43546
rect 14382 43494 14394 43546
rect 14394 43494 14408 43546
rect 14432 43494 14446 43546
rect 14446 43494 14458 43546
rect 14458 43494 14488 43546
rect 14512 43494 14522 43546
rect 14522 43494 14568 43546
rect 14272 43492 14328 43494
rect 14352 43492 14408 43494
rect 14432 43492 14488 43494
rect 14512 43492 14568 43494
rect 18711 43546 18767 43548
rect 18791 43546 18847 43548
rect 18871 43546 18927 43548
rect 18951 43546 19007 43548
rect 18711 43494 18757 43546
rect 18757 43494 18767 43546
rect 18791 43494 18821 43546
rect 18821 43494 18833 43546
rect 18833 43494 18847 43546
rect 18871 43494 18885 43546
rect 18885 43494 18897 43546
rect 18897 43494 18927 43546
rect 18951 43494 18961 43546
rect 18961 43494 19007 43546
rect 18711 43492 18767 43494
rect 18791 43492 18847 43494
rect 18871 43492 18927 43494
rect 18951 43492 19007 43494
rect 3175 43002 3231 43004
rect 3255 43002 3311 43004
rect 3335 43002 3391 43004
rect 3415 43002 3471 43004
rect 3175 42950 3221 43002
rect 3221 42950 3231 43002
rect 3255 42950 3285 43002
rect 3285 42950 3297 43002
rect 3297 42950 3311 43002
rect 3335 42950 3349 43002
rect 3349 42950 3361 43002
rect 3361 42950 3391 43002
rect 3415 42950 3425 43002
rect 3425 42950 3471 43002
rect 3175 42948 3231 42950
rect 3255 42948 3311 42950
rect 3335 42948 3391 42950
rect 3415 42948 3471 42950
rect 7614 43002 7670 43004
rect 7694 43002 7750 43004
rect 7774 43002 7830 43004
rect 7854 43002 7910 43004
rect 7614 42950 7660 43002
rect 7660 42950 7670 43002
rect 7694 42950 7724 43002
rect 7724 42950 7736 43002
rect 7736 42950 7750 43002
rect 7774 42950 7788 43002
rect 7788 42950 7800 43002
rect 7800 42950 7830 43002
rect 7854 42950 7864 43002
rect 7864 42950 7910 43002
rect 7614 42948 7670 42950
rect 7694 42948 7750 42950
rect 7774 42948 7830 42950
rect 7854 42948 7910 42950
rect 12053 43002 12109 43004
rect 12133 43002 12189 43004
rect 12213 43002 12269 43004
rect 12293 43002 12349 43004
rect 12053 42950 12099 43002
rect 12099 42950 12109 43002
rect 12133 42950 12163 43002
rect 12163 42950 12175 43002
rect 12175 42950 12189 43002
rect 12213 42950 12227 43002
rect 12227 42950 12239 43002
rect 12239 42950 12269 43002
rect 12293 42950 12303 43002
rect 12303 42950 12349 43002
rect 12053 42948 12109 42950
rect 12133 42948 12189 42950
rect 12213 42948 12269 42950
rect 12293 42948 12349 42950
rect 16492 43002 16548 43004
rect 16572 43002 16628 43004
rect 16652 43002 16708 43004
rect 16732 43002 16788 43004
rect 16492 42950 16538 43002
rect 16538 42950 16548 43002
rect 16572 42950 16602 43002
rect 16602 42950 16614 43002
rect 16614 42950 16628 43002
rect 16652 42950 16666 43002
rect 16666 42950 16678 43002
rect 16678 42950 16708 43002
rect 16732 42950 16742 43002
rect 16742 42950 16788 43002
rect 16492 42948 16548 42950
rect 16572 42948 16628 42950
rect 16652 42948 16708 42950
rect 16732 42948 16788 42950
rect 5394 42458 5450 42460
rect 5474 42458 5530 42460
rect 5554 42458 5610 42460
rect 5634 42458 5690 42460
rect 5394 42406 5440 42458
rect 5440 42406 5450 42458
rect 5474 42406 5504 42458
rect 5504 42406 5516 42458
rect 5516 42406 5530 42458
rect 5554 42406 5568 42458
rect 5568 42406 5580 42458
rect 5580 42406 5610 42458
rect 5634 42406 5644 42458
rect 5644 42406 5690 42458
rect 5394 42404 5450 42406
rect 5474 42404 5530 42406
rect 5554 42404 5610 42406
rect 5634 42404 5690 42406
rect 9833 42458 9889 42460
rect 9913 42458 9969 42460
rect 9993 42458 10049 42460
rect 10073 42458 10129 42460
rect 9833 42406 9879 42458
rect 9879 42406 9889 42458
rect 9913 42406 9943 42458
rect 9943 42406 9955 42458
rect 9955 42406 9969 42458
rect 9993 42406 10007 42458
rect 10007 42406 10019 42458
rect 10019 42406 10049 42458
rect 10073 42406 10083 42458
rect 10083 42406 10129 42458
rect 9833 42404 9889 42406
rect 9913 42404 9969 42406
rect 9993 42404 10049 42406
rect 10073 42404 10129 42406
rect 14272 42458 14328 42460
rect 14352 42458 14408 42460
rect 14432 42458 14488 42460
rect 14512 42458 14568 42460
rect 14272 42406 14318 42458
rect 14318 42406 14328 42458
rect 14352 42406 14382 42458
rect 14382 42406 14394 42458
rect 14394 42406 14408 42458
rect 14432 42406 14446 42458
rect 14446 42406 14458 42458
rect 14458 42406 14488 42458
rect 14512 42406 14522 42458
rect 14522 42406 14568 42458
rect 14272 42404 14328 42406
rect 14352 42404 14408 42406
rect 14432 42404 14488 42406
rect 14512 42404 14568 42406
rect 18711 42458 18767 42460
rect 18791 42458 18847 42460
rect 18871 42458 18927 42460
rect 18951 42458 19007 42460
rect 18711 42406 18757 42458
rect 18757 42406 18767 42458
rect 18791 42406 18821 42458
rect 18821 42406 18833 42458
rect 18833 42406 18847 42458
rect 18871 42406 18885 42458
rect 18885 42406 18897 42458
rect 18897 42406 18927 42458
rect 18951 42406 18961 42458
rect 18961 42406 19007 42458
rect 18711 42404 18767 42406
rect 18791 42404 18847 42406
rect 18871 42404 18927 42406
rect 18951 42404 19007 42406
rect 3175 41914 3231 41916
rect 3255 41914 3311 41916
rect 3335 41914 3391 41916
rect 3415 41914 3471 41916
rect 3175 41862 3221 41914
rect 3221 41862 3231 41914
rect 3255 41862 3285 41914
rect 3285 41862 3297 41914
rect 3297 41862 3311 41914
rect 3335 41862 3349 41914
rect 3349 41862 3361 41914
rect 3361 41862 3391 41914
rect 3415 41862 3425 41914
rect 3425 41862 3471 41914
rect 3175 41860 3231 41862
rect 3255 41860 3311 41862
rect 3335 41860 3391 41862
rect 3415 41860 3471 41862
rect 7614 41914 7670 41916
rect 7694 41914 7750 41916
rect 7774 41914 7830 41916
rect 7854 41914 7910 41916
rect 7614 41862 7660 41914
rect 7660 41862 7670 41914
rect 7694 41862 7724 41914
rect 7724 41862 7736 41914
rect 7736 41862 7750 41914
rect 7774 41862 7788 41914
rect 7788 41862 7800 41914
rect 7800 41862 7830 41914
rect 7854 41862 7864 41914
rect 7864 41862 7910 41914
rect 7614 41860 7670 41862
rect 7694 41860 7750 41862
rect 7774 41860 7830 41862
rect 7854 41860 7910 41862
rect 12053 41914 12109 41916
rect 12133 41914 12189 41916
rect 12213 41914 12269 41916
rect 12293 41914 12349 41916
rect 12053 41862 12099 41914
rect 12099 41862 12109 41914
rect 12133 41862 12163 41914
rect 12163 41862 12175 41914
rect 12175 41862 12189 41914
rect 12213 41862 12227 41914
rect 12227 41862 12239 41914
rect 12239 41862 12269 41914
rect 12293 41862 12303 41914
rect 12303 41862 12349 41914
rect 12053 41860 12109 41862
rect 12133 41860 12189 41862
rect 12213 41860 12269 41862
rect 12293 41860 12349 41862
rect 16492 41914 16548 41916
rect 16572 41914 16628 41916
rect 16652 41914 16708 41916
rect 16732 41914 16788 41916
rect 16492 41862 16538 41914
rect 16538 41862 16548 41914
rect 16572 41862 16602 41914
rect 16602 41862 16614 41914
rect 16614 41862 16628 41914
rect 16652 41862 16666 41914
rect 16666 41862 16678 41914
rect 16678 41862 16708 41914
rect 16732 41862 16742 41914
rect 16742 41862 16788 41914
rect 16492 41860 16548 41862
rect 16572 41860 16628 41862
rect 16652 41860 16708 41862
rect 16732 41860 16788 41862
rect 5394 41370 5450 41372
rect 5474 41370 5530 41372
rect 5554 41370 5610 41372
rect 5634 41370 5690 41372
rect 5394 41318 5440 41370
rect 5440 41318 5450 41370
rect 5474 41318 5504 41370
rect 5504 41318 5516 41370
rect 5516 41318 5530 41370
rect 5554 41318 5568 41370
rect 5568 41318 5580 41370
rect 5580 41318 5610 41370
rect 5634 41318 5644 41370
rect 5644 41318 5690 41370
rect 5394 41316 5450 41318
rect 5474 41316 5530 41318
rect 5554 41316 5610 41318
rect 5634 41316 5690 41318
rect 9833 41370 9889 41372
rect 9913 41370 9969 41372
rect 9993 41370 10049 41372
rect 10073 41370 10129 41372
rect 9833 41318 9879 41370
rect 9879 41318 9889 41370
rect 9913 41318 9943 41370
rect 9943 41318 9955 41370
rect 9955 41318 9969 41370
rect 9993 41318 10007 41370
rect 10007 41318 10019 41370
rect 10019 41318 10049 41370
rect 10073 41318 10083 41370
rect 10083 41318 10129 41370
rect 9833 41316 9889 41318
rect 9913 41316 9969 41318
rect 9993 41316 10049 41318
rect 10073 41316 10129 41318
rect 14272 41370 14328 41372
rect 14352 41370 14408 41372
rect 14432 41370 14488 41372
rect 14512 41370 14568 41372
rect 14272 41318 14318 41370
rect 14318 41318 14328 41370
rect 14352 41318 14382 41370
rect 14382 41318 14394 41370
rect 14394 41318 14408 41370
rect 14432 41318 14446 41370
rect 14446 41318 14458 41370
rect 14458 41318 14488 41370
rect 14512 41318 14522 41370
rect 14522 41318 14568 41370
rect 14272 41316 14328 41318
rect 14352 41316 14408 41318
rect 14432 41316 14488 41318
rect 14512 41316 14568 41318
rect 18711 41370 18767 41372
rect 18791 41370 18847 41372
rect 18871 41370 18927 41372
rect 18951 41370 19007 41372
rect 18711 41318 18757 41370
rect 18757 41318 18767 41370
rect 18791 41318 18821 41370
rect 18821 41318 18833 41370
rect 18833 41318 18847 41370
rect 18871 41318 18885 41370
rect 18885 41318 18897 41370
rect 18897 41318 18927 41370
rect 18951 41318 18961 41370
rect 18961 41318 19007 41370
rect 18711 41316 18767 41318
rect 18791 41316 18847 41318
rect 18871 41316 18927 41318
rect 18951 41316 19007 41318
rect 938 9016 994 9072
rect 938 5480 994 5536
rect 1766 26560 1822 26616
rect 2042 19372 2098 19408
rect 3175 40826 3231 40828
rect 3255 40826 3311 40828
rect 3335 40826 3391 40828
rect 3415 40826 3471 40828
rect 3175 40774 3221 40826
rect 3221 40774 3231 40826
rect 3255 40774 3285 40826
rect 3285 40774 3297 40826
rect 3297 40774 3311 40826
rect 3335 40774 3349 40826
rect 3349 40774 3361 40826
rect 3361 40774 3391 40826
rect 3415 40774 3425 40826
rect 3425 40774 3471 40826
rect 3175 40772 3231 40774
rect 3255 40772 3311 40774
rect 3335 40772 3391 40774
rect 3415 40772 3471 40774
rect 7614 40826 7670 40828
rect 7694 40826 7750 40828
rect 7774 40826 7830 40828
rect 7854 40826 7910 40828
rect 7614 40774 7660 40826
rect 7660 40774 7670 40826
rect 7694 40774 7724 40826
rect 7724 40774 7736 40826
rect 7736 40774 7750 40826
rect 7774 40774 7788 40826
rect 7788 40774 7800 40826
rect 7800 40774 7830 40826
rect 7854 40774 7864 40826
rect 7864 40774 7910 40826
rect 7614 40772 7670 40774
rect 7694 40772 7750 40774
rect 7774 40772 7830 40774
rect 7854 40772 7910 40774
rect 12053 40826 12109 40828
rect 12133 40826 12189 40828
rect 12213 40826 12269 40828
rect 12293 40826 12349 40828
rect 12053 40774 12099 40826
rect 12099 40774 12109 40826
rect 12133 40774 12163 40826
rect 12163 40774 12175 40826
rect 12175 40774 12189 40826
rect 12213 40774 12227 40826
rect 12227 40774 12239 40826
rect 12239 40774 12269 40826
rect 12293 40774 12303 40826
rect 12303 40774 12349 40826
rect 12053 40772 12109 40774
rect 12133 40772 12189 40774
rect 12213 40772 12269 40774
rect 12293 40772 12349 40774
rect 16492 40826 16548 40828
rect 16572 40826 16628 40828
rect 16652 40826 16708 40828
rect 16732 40826 16788 40828
rect 16492 40774 16538 40826
rect 16538 40774 16548 40826
rect 16572 40774 16602 40826
rect 16602 40774 16614 40826
rect 16614 40774 16628 40826
rect 16652 40774 16666 40826
rect 16666 40774 16678 40826
rect 16678 40774 16708 40826
rect 16732 40774 16742 40826
rect 16742 40774 16788 40826
rect 16492 40772 16548 40774
rect 16572 40772 16628 40774
rect 16652 40772 16708 40774
rect 16732 40772 16788 40774
rect 5394 40282 5450 40284
rect 5474 40282 5530 40284
rect 5554 40282 5610 40284
rect 5634 40282 5690 40284
rect 5394 40230 5440 40282
rect 5440 40230 5450 40282
rect 5474 40230 5504 40282
rect 5504 40230 5516 40282
rect 5516 40230 5530 40282
rect 5554 40230 5568 40282
rect 5568 40230 5580 40282
rect 5580 40230 5610 40282
rect 5634 40230 5644 40282
rect 5644 40230 5690 40282
rect 5394 40228 5450 40230
rect 5474 40228 5530 40230
rect 5554 40228 5610 40230
rect 5634 40228 5690 40230
rect 9833 40282 9889 40284
rect 9913 40282 9969 40284
rect 9993 40282 10049 40284
rect 10073 40282 10129 40284
rect 9833 40230 9879 40282
rect 9879 40230 9889 40282
rect 9913 40230 9943 40282
rect 9943 40230 9955 40282
rect 9955 40230 9969 40282
rect 9993 40230 10007 40282
rect 10007 40230 10019 40282
rect 10019 40230 10049 40282
rect 10073 40230 10083 40282
rect 10083 40230 10129 40282
rect 9833 40228 9889 40230
rect 9913 40228 9969 40230
rect 9993 40228 10049 40230
rect 10073 40228 10129 40230
rect 14272 40282 14328 40284
rect 14352 40282 14408 40284
rect 14432 40282 14488 40284
rect 14512 40282 14568 40284
rect 14272 40230 14318 40282
rect 14318 40230 14328 40282
rect 14352 40230 14382 40282
rect 14382 40230 14394 40282
rect 14394 40230 14408 40282
rect 14432 40230 14446 40282
rect 14446 40230 14458 40282
rect 14458 40230 14488 40282
rect 14512 40230 14522 40282
rect 14522 40230 14568 40282
rect 14272 40228 14328 40230
rect 14352 40228 14408 40230
rect 14432 40228 14488 40230
rect 14512 40228 14568 40230
rect 18711 40282 18767 40284
rect 18791 40282 18847 40284
rect 18871 40282 18927 40284
rect 18951 40282 19007 40284
rect 18711 40230 18757 40282
rect 18757 40230 18767 40282
rect 18791 40230 18821 40282
rect 18821 40230 18833 40282
rect 18833 40230 18847 40282
rect 18871 40230 18885 40282
rect 18885 40230 18897 40282
rect 18897 40230 18927 40282
rect 18951 40230 18961 40282
rect 18961 40230 19007 40282
rect 18711 40228 18767 40230
rect 18791 40228 18847 40230
rect 18871 40228 18927 40230
rect 18951 40228 19007 40230
rect 3175 39738 3231 39740
rect 3255 39738 3311 39740
rect 3335 39738 3391 39740
rect 3415 39738 3471 39740
rect 3175 39686 3221 39738
rect 3221 39686 3231 39738
rect 3255 39686 3285 39738
rect 3285 39686 3297 39738
rect 3297 39686 3311 39738
rect 3335 39686 3349 39738
rect 3349 39686 3361 39738
rect 3361 39686 3391 39738
rect 3415 39686 3425 39738
rect 3425 39686 3471 39738
rect 3175 39684 3231 39686
rect 3255 39684 3311 39686
rect 3335 39684 3391 39686
rect 3415 39684 3471 39686
rect 7614 39738 7670 39740
rect 7694 39738 7750 39740
rect 7774 39738 7830 39740
rect 7854 39738 7910 39740
rect 7614 39686 7660 39738
rect 7660 39686 7670 39738
rect 7694 39686 7724 39738
rect 7724 39686 7736 39738
rect 7736 39686 7750 39738
rect 7774 39686 7788 39738
rect 7788 39686 7800 39738
rect 7800 39686 7830 39738
rect 7854 39686 7864 39738
rect 7864 39686 7910 39738
rect 7614 39684 7670 39686
rect 7694 39684 7750 39686
rect 7774 39684 7830 39686
rect 7854 39684 7910 39686
rect 12053 39738 12109 39740
rect 12133 39738 12189 39740
rect 12213 39738 12269 39740
rect 12293 39738 12349 39740
rect 12053 39686 12099 39738
rect 12099 39686 12109 39738
rect 12133 39686 12163 39738
rect 12163 39686 12175 39738
rect 12175 39686 12189 39738
rect 12213 39686 12227 39738
rect 12227 39686 12239 39738
rect 12239 39686 12269 39738
rect 12293 39686 12303 39738
rect 12303 39686 12349 39738
rect 12053 39684 12109 39686
rect 12133 39684 12189 39686
rect 12213 39684 12269 39686
rect 12293 39684 12349 39686
rect 16492 39738 16548 39740
rect 16572 39738 16628 39740
rect 16652 39738 16708 39740
rect 16732 39738 16788 39740
rect 16492 39686 16538 39738
rect 16538 39686 16548 39738
rect 16572 39686 16602 39738
rect 16602 39686 16614 39738
rect 16614 39686 16628 39738
rect 16652 39686 16666 39738
rect 16666 39686 16678 39738
rect 16678 39686 16708 39738
rect 16732 39686 16742 39738
rect 16742 39686 16788 39738
rect 16492 39684 16548 39686
rect 16572 39684 16628 39686
rect 16652 39684 16708 39686
rect 16732 39684 16788 39686
rect 5394 39194 5450 39196
rect 5474 39194 5530 39196
rect 5554 39194 5610 39196
rect 5634 39194 5690 39196
rect 5394 39142 5440 39194
rect 5440 39142 5450 39194
rect 5474 39142 5504 39194
rect 5504 39142 5516 39194
rect 5516 39142 5530 39194
rect 5554 39142 5568 39194
rect 5568 39142 5580 39194
rect 5580 39142 5610 39194
rect 5634 39142 5644 39194
rect 5644 39142 5690 39194
rect 5394 39140 5450 39142
rect 5474 39140 5530 39142
rect 5554 39140 5610 39142
rect 5634 39140 5690 39142
rect 9833 39194 9889 39196
rect 9913 39194 9969 39196
rect 9993 39194 10049 39196
rect 10073 39194 10129 39196
rect 9833 39142 9879 39194
rect 9879 39142 9889 39194
rect 9913 39142 9943 39194
rect 9943 39142 9955 39194
rect 9955 39142 9969 39194
rect 9993 39142 10007 39194
rect 10007 39142 10019 39194
rect 10019 39142 10049 39194
rect 10073 39142 10083 39194
rect 10083 39142 10129 39194
rect 9833 39140 9889 39142
rect 9913 39140 9969 39142
rect 9993 39140 10049 39142
rect 10073 39140 10129 39142
rect 14272 39194 14328 39196
rect 14352 39194 14408 39196
rect 14432 39194 14488 39196
rect 14512 39194 14568 39196
rect 14272 39142 14318 39194
rect 14318 39142 14328 39194
rect 14352 39142 14382 39194
rect 14382 39142 14394 39194
rect 14394 39142 14408 39194
rect 14432 39142 14446 39194
rect 14446 39142 14458 39194
rect 14458 39142 14488 39194
rect 14512 39142 14522 39194
rect 14522 39142 14568 39194
rect 14272 39140 14328 39142
rect 14352 39140 14408 39142
rect 14432 39140 14488 39142
rect 14512 39140 14568 39142
rect 18711 39194 18767 39196
rect 18791 39194 18847 39196
rect 18871 39194 18927 39196
rect 18951 39194 19007 39196
rect 18711 39142 18757 39194
rect 18757 39142 18767 39194
rect 18791 39142 18821 39194
rect 18821 39142 18833 39194
rect 18833 39142 18847 39194
rect 18871 39142 18885 39194
rect 18885 39142 18897 39194
rect 18897 39142 18927 39194
rect 18951 39142 18961 39194
rect 18961 39142 19007 39194
rect 18711 39140 18767 39142
rect 18791 39140 18847 39142
rect 18871 39140 18927 39142
rect 18951 39140 19007 39142
rect 3175 38650 3231 38652
rect 3255 38650 3311 38652
rect 3335 38650 3391 38652
rect 3415 38650 3471 38652
rect 3175 38598 3221 38650
rect 3221 38598 3231 38650
rect 3255 38598 3285 38650
rect 3285 38598 3297 38650
rect 3297 38598 3311 38650
rect 3335 38598 3349 38650
rect 3349 38598 3361 38650
rect 3361 38598 3391 38650
rect 3415 38598 3425 38650
rect 3425 38598 3471 38650
rect 3175 38596 3231 38598
rect 3255 38596 3311 38598
rect 3335 38596 3391 38598
rect 3415 38596 3471 38598
rect 7614 38650 7670 38652
rect 7694 38650 7750 38652
rect 7774 38650 7830 38652
rect 7854 38650 7910 38652
rect 7614 38598 7660 38650
rect 7660 38598 7670 38650
rect 7694 38598 7724 38650
rect 7724 38598 7736 38650
rect 7736 38598 7750 38650
rect 7774 38598 7788 38650
rect 7788 38598 7800 38650
rect 7800 38598 7830 38650
rect 7854 38598 7864 38650
rect 7864 38598 7910 38650
rect 7614 38596 7670 38598
rect 7694 38596 7750 38598
rect 7774 38596 7830 38598
rect 7854 38596 7910 38598
rect 12053 38650 12109 38652
rect 12133 38650 12189 38652
rect 12213 38650 12269 38652
rect 12293 38650 12349 38652
rect 12053 38598 12099 38650
rect 12099 38598 12109 38650
rect 12133 38598 12163 38650
rect 12163 38598 12175 38650
rect 12175 38598 12189 38650
rect 12213 38598 12227 38650
rect 12227 38598 12239 38650
rect 12239 38598 12269 38650
rect 12293 38598 12303 38650
rect 12303 38598 12349 38650
rect 12053 38596 12109 38598
rect 12133 38596 12189 38598
rect 12213 38596 12269 38598
rect 12293 38596 12349 38598
rect 16492 38650 16548 38652
rect 16572 38650 16628 38652
rect 16652 38650 16708 38652
rect 16732 38650 16788 38652
rect 16492 38598 16538 38650
rect 16538 38598 16548 38650
rect 16572 38598 16602 38650
rect 16602 38598 16614 38650
rect 16614 38598 16628 38650
rect 16652 38598 16666 38650
rect 16666 38598 16678 38650
rect 16678 38598 16708 38650
rect 16732 38598 16742 38650
rect 16742 38598 16788 38650
rect 16492 38596 16548 38598
rect 16572 38596 16628 38598
rect 16652 38596 16708 38598
rect 16732 38596 16788 38598
rect 5394 38106 5450 38108
rect 5474 38106 5530 38108
rect 5554 38106 5610 38108
rect 5634 38106 5690 38108
rect 5394 38054 5440 38106
rect 5440 38054 5450 38106
rect 5474 38054 5504 38106
rect 5504 38054 5516 38106
rect 5516 38054 5530 38106
rect 5554 38054 5568 38106
rect 5568 38054 5580 38106
rect 5580 38054 5610 38106
rect 5634 38054 5644 38106
rect 5644 38054 5690 38106
rect 5394 38052 5450 38054
rect 5474 38052 5530 38054
rect 5554 38052 5610 38054
rect 5634 38052 5690 38054
rect 9833 38106 9889 38108
rect 9913 38106 9969 38108
rect 9993 38106 10049 38108
rect 10073 38106 10129 38108
rect 9833 38054 9879 38106
rect 9879 38054 9889 38106
rect 9913 38054 9943 38106
rect 9943 38054 9955 38106
rect 9955 38054 9969 38106
rect 9993 38054 10007 38106
rect 10007 38054 10019 38106
rect 10019 38054 10049 38106
rect 10073 38054 10083 38106
rect 10083 38054 10129 38106
rect 9833 38052 9889 38054
rect 9913 38052 9969 38054
rect 9993 38052 10049 38054
rect 10073 38052 10129 38054
rect 14272 38106 14328 38108
rect 14352 38106 14408 38108
rect 14432 38106 14488 38108
rect 14512 38106 14568 38108
rect 14272 38054 14318 38106
rect 14318 38054 14328 38106
rect 14352 38054 14382 38106
rect 14382 38054 14394 38106
rect 14394 38054 14408 38106
rect 14432 38054 14446 38106
rect 14446 38054 14458 38106
rect 14458 38054 14488 38106
rect 14512 38054 14522 38106
rect 14522 38054 14568 38106
rect 14272 38052 14328 38054
rect 14352 38052 14408 38054
rect 14432 38052 14488 38054
rect 14512 38052 14568 38054
rect 18711 38106 18767 38108
rect 18791 38106 18847 38108
rect 18871 38106 18927 38108
rect 18951 38106 19007 38108
rect 18711 38054 18757 38106
rect 18757 38054 18767 38106
rect 18791 38054 18821 38106
rect 18821 38054 18833 38106
rect 18833 38054 18847 38106
rect 18871 38054 18885 38106
rect 18885 38054 18897 38106
rect 18897 38054 18927 38106
rect 18951 38054 18961 38106
rect 18961 38054 19007 38106
rect 18711 38052 18767 38054
rect 18791 38052 18847 38054
rect 18871 38052 18927 38054
rect 18951 38052 19007 38054
rect 3175 37562 3231 37564
rect 3255 37562 3311 37564
rect 3335 37562 3391 37564
rect 3415 37562 3471 37564
rect 3175 37510 3221 37562
rect 3221 37510 3231 37562
rect 3255 37510 3285 37562
rect 3285 37510 3297 37562
rect 3297 37510 3311 37562
rect 3335 37510 3349 37562
rect 3349 37510 3361 37562
rect 3361 37510 3391 37562
rect 3415 37510 3425 37562
rect 3425 37510 3471 37562
rect 3175 37508 3231 37510
rect 3255 37508 3311 37510
rect 3335 37508 3391 37510
rect 3415 37508 3471 37510
rect 7614 37562 7670 37564
rect 7694 37562 7750 37564
rect 7774 37562 7830 37564
rect 7854 37562 7910 37564
rect 7614 37510 7660 37562
rect 7660 37510 7670 37562
rect 7694 37510 7724 37562
rect 7724 37510 7736 37562
rect 7736 37510 7750 37562
rect 7774 37510 7788 37562
rect 7788 37510 7800 37562
rect 7800 37510 7830 37562
rect 7854 37510 7864 37562
rect 7864 37510 7910 37562
rect 7614 37508 7670 37510
rect 7694 37508 7750 37510
rect 7774 37508 7830 37510
rect 7854 37508 7910 37510
rect 12053 37562 12109 37564
rect 12133 37562 12189 37564
rect 12213 37562 12269 37564
rect 12293 37562 12349 37564
rect 12053 37510 12099 37562
rect 12099 37510 12109 37562
rect 12133 37510 12163 37562
rect 12163 37510 12175 37562
rect 12175 37510 12189 37562
rect 12213 37510 12227 37562
rect 12227 37510 12239 37562
rect 12239 37510 12269 37562
rect 12293 37510 12303 37562
rect 12303 37510 12349 37562
rect 12053 37508 12109 37510
rect 12133 37508 12189 37510
rect 12213 37508 12269 37510
rect 12293 37508 12349 37510
rect 16492 37562 16548 37564
rect 16572 37562 16628 37564
rect 16652 37562 16708 37564
rect 16732 37562 16788 37564
rect 16492 37510 16538 37562
rect 16538 37510 16548 37562
rect 16572 37510 16602 37562
rect 16602 37510 16614 37562
rect 16614 37510 16628 37562
rect 16652 37510 16666 37562
rect 16666 37510 16678 37562
rect 16678 37510 16708 37562
rect 16732 37510 16742 37562
rect 16742 37510 16788 37562
rect 16492 37508 16548 37510
rect 16572 37508 16628 37510
rect 16652 37508 16708 37510
rect 16732 37508 16788 37510
rect 5394 37018 5450 37020
rect 5474 37018 5530 37020
rect 5554 37018 5610 37020
rect 5634 37018 5690 37020
rect 5394 36966 5440 37018
rect 5440 36966 5450 37018
rect 5474 36966 5504 37018
rect 5504 36966 5516 37018
rect 5516 36966 5530 37018
rect 5554 36966 5568 37018
rect 5568 36966 5580 37018
rect 5580 36966 5610 37018
rect 5634 36966 5644 37018
rect 5644 36966 5690 37018
rect 5394 36964 5450 36966
rect 5474 36964 5530 36966
rect 5554 36964 5610 36966
rect 5634 36964 5690 36966
rect 9833 37018 9889 37020
rect 9913 37018 9969 37020
rect 9993 37018 10049 37020
rect 10073 37018 10129 37020
rect 9833 36966 9879 37018
rect 9879 36966 9889 37018
rect 9913 36966 9943 37018
rect 9943 36966 9955 37018
rect 9955 36966 9969 37018
rect 9993 36966 10007 37018
rect 10007 36966 10019 37018
rect 10019 36966 10049 37018
rect 10073 36966 10083 37018
rect 10083 36966 10129 37018
rect 9833 36964 9889 36966
rect 9913 36964 9969 36966
rect 9993 36964 10049 36966
rect 10073 36964 10129 36966
rect 14272 37018 14328 37020
rect 14352 37018 14408 37020
rect 14432 37018 14488 37020
rect 14512 37018 14568 37020
rect 14272 36966 14318 37018
rect 14318 36966 14328 37018
rect 14352 36966 14382 37018
rect 14382 36966 14394 37018
rect 14394 36966 14408 37018
rect 14432 36966 14446 37018
rect 14446 36966 14458 37018
rect 14458 36966 14488 37018
rect 14512 36966 14522 37018
rect 14522 36966 14568 37018
rect 14272 36964 14328 36966
rect 14352 36964 14408 36966
rect 14432 36964 14488 36966
rect 14512 36964 14568 36966
rect 18711 37018 18767 37020
rect 18791 37018 18847 37020
rect 18871 37018 18927 37020
rect 18951 37018 19007 37020
rect 18711 36966 18757 37018
rect 18757 36966 18767 37018
rect 18791 36966 18821 37018
rect 18821 36966 18833 37018
rect 18833 36966 18847 37018
rect 18871 36966 18885 37018
rect 18885 36966 18897 37018
rect 18897 36966 18927 37018
rect 18951 36966 18961 37018
rect 18961 36966 19007 37018
rect 18711 36964 18767 36966
rect 18791 36964 18847 36966
rect 18871 36964 18927 36966
rect 18951 36964 19007 36966
rect 3175 36474 3231 36476
rect 3255 36474 3311 36476
rect 3335 36474 3391 36476
rect 3415 36474 3471 36476
rect 3175 36422 3221 36474
rect 3221 36422 3231 36474
rect 3255 36422 3285 36474
rect 3285 36422 3297 36474
rect 3297 36422 3311 36474
rect 3335 36422 3349 36474
rect 3349 36422 3361 36474
rect 3361 36422 3391 36474
rect 3415 36422 3425 36474
rect 3425 36422 3471 36474
rect 3175 36420 3231 36422
rect 3255 36420 3311 36422
rect 3335 36420 3391 36422
rect 3415 36420 3471 36422
rect 7614 36474 7670 36476
rect 7694 36474 7750 36476
rect 7774 36474 7830 36476
rect 7854 36474 7910 36476
rect 7614 36422 7660 36474
rect 7660 36422 7670 36474
rect 7694 36422 7724 36474
rect 7724 36422 7736 36474
rect 7736 36422 7750 36474
rect 7774 36422 7788 36474
rect 7788 36422 7800 36474
rect 7800 36422 7830 36474
rect 7854 36422 7864 36474
rect 7864 36422 7910 36474
rect 7614 36420 7670 36422
rect 7694 36420 7750 36422
rect 7774 36420 7830 36422
rect 7854 36420 7910 36422
rect 12053 36474 12109 36476
rect 12133 36474 12189 36476
rect 12213 36474 12269 36476
rect 12293 36474 12349 36476
rect 12053 36422 12099 36474
rect 12099 36422 12109 36474
rect 12133 36422 12163 36474
rect 12163 36422 12175 36474
rect 12175 36422 12189 36474
rect 12213 36422 12227 36474
rect 12227 36422 12239 36474
rect 12239 36422 12269 36474
rect 12293 36422 12303 36474
rect 12303 36422 12349 36474
rect 12053 36420 12109 36422
rect 12133 36420 12189 36422
rect 12213 36420 12269 36422
rect 12293 36420 12349 36422
rect 16492 36474 16548 36476
rect 16572 36474 16628 36476
rect 16652 36474 16708 36476
rect 16732 36474 16788 36476
rect 16492 36422 16538 36474
rect 16538 36422 16548 36474
rect 16572 36422 16602 36474
rect 16602 36422 16614 36474
rect 16614 36422 16628 36474
rect 16652 36422 16666 36474
rect 16666 36422 16678 36474
rect 16678 36422 16708 36474
rect 16732 36422 16742 36474
rect 16742 36422 16788 36474
rect 16492 36420 16548 36422
rect 16572 36420 16628 36422
rect 16652 36420 16708 36422
rect 16732 36420 16788 36422
rect 5394 35930 5450 35932
rect 5474 35930 5530 35932
rect 5554 35930 5610 35932
rect 5634 35930 5690 35932
rect 5394 35878 5440 35930
rect 5440 35878 5450 35930
rect 5474 35878 5504 35930
rect 5504 35878 5516 35930
rect 5516 35878 5530 35930
rect 5554 35878 5568 35930
rect 5568 35878 5580 35930
rect 5580 35878 5610 35930
rect 5634 35878 5644 35930
rect 5644 35878 5690 35930
rect 5394 35876 5450 35878
rect 5474 35876 5530 35878
rect 5554 35876 5610 35878
rect 5634 35876 5690 35878
rect 3175 35386 3231 35388
rect 3255 35386 3311 35388
rect 3335 35386 3391 35388
rect 3415 35386 3471 35388
rect 3175 35334 3221 35386
rect 3221 35334 3231 35386
rect 3255 35334 3285 35386
rect 3285 35334 3297 35386
rect 3297 35334 3311 35386
rect 3335 35334 3349 35386
rect 3349 35334 3361 35386
rect 3361 35334 3391 35386
rect 3415 35334 3425 35386
rect 3425 35334 3471 35386
rect 3175 35332 3231 35334
rect 3255 35332 3311 35334
rect 3335 35332 3391 35334
rect 3415 35332 3471 35334
rect 3175 34298 3231 34300
rect 3255 34298 3311 34300
rect 3335 34298 3391 34300
rect 3415 34298 3471 34300
rect 3175 34246 3221 34298
rect 3221 34246 3231 34298
rect 3255 34246 3285 34298
rect 3285 34246 3297 34298
rect 3297 34246 3311 34298
rect 3335 34246 3349 34298
rect 3349 34246 3361 34298
rect 3361 34246 3391 34298
rect 3415 34246 3425 34298
rect 3425 34246 3471 34298
rect 3175 34244 3231 34246
rect 3255 34244 3311 34246
rect 3335 34244 3391 34246
rect 3415 34244 3471 34246
rect 3175 33210 3231 33212
rect 3255 33210 3311 33212
rect 3335 33210 3391 33212
rect 3415 33210 3471 33212
rect 3175 33158 3221 33210
rect 3221 33158 3231 33210
rect 3255 33158 3285 33210
rect 3285 33158 3297 33210
rect 3297 33158 3311 33210
rect 3335 33158 3349 33210
rect 3349 33158 3361 33210
rect 3361 33158 3391 33210
rect 3415 33158 3425 33210
rect 3425 33158 3471 33210
rect 3175 33156 3231 33158
rect 3255 33156 3311 33158
rect 3335 33156 3391 33158
rect 3415 33156 3471 33158
rect 3175 32122 3231 32124
rect 3255 32122 3311 32124
rect 3335 32122 3391 32124
rect 3415 32122 3471 32124
rect 3175 32070 3221 32122
rect 3221 32070 3231 32122
rect 3255 32070 3285 32122
rect 3285 32070 3297 32122
rect 3297 32070 3311 32122
rect 3335 32070 3349 32122
rect 3349 32070 3361 32122
rect 3361 32070 3391 32122
rect 3415 32070 3425 32122
rect 3425 32070 3471 32122
rect 3175 32068 3231 32070
rect 3255 32068 3311 32070
rect 3335 32068 3391 32070
rect 3415 32068 3471 32070
rect 3175 31034 3231 31036
rect 3255 31034 3311 31036
rect 3335 31034 3391 31036
rect 3415 31034 3471 31036
rect 3175 30982 3221 31034
rect 3221 30982 3231 31034
rect 3255 30982 3285 31034
rect 3285 30982 3297 31034
rect 3297 30982 3311 31034
rect 3335 30982 3349 31034
rect 3349 30982 3361 31034
rect 3361 30982 3391 31034
rect 3415 30982 3425 31034
rect 3425 30982 3471 31034
rect 3175 30980 3231 30982
rect 3255 30980 3311 30982
rect 3335 30980 3391 30982
rect 3415 30980 3471 30982
rect 5394 34842 5450 34844
rect 5474 34842 5530 34844
rect 5554 34842 5610 34844
rect 5634 34842 5690 34844
rect 5394 34790 5440 34842
rect 5440 34790 5450 34842
rect 5474 34790 5504 34842
rect 5504 34790 5516 34842
rect 5516 34790 5530 34842
rect 5554 34790 5568 34842
rect 5568 34790 5580 34842
rect 5580 34790 5610 34842
rect 5634 34790 5644 34842
rect 5644 34790 5690 34842
rect 5394 34788 5450 34790
rect 5474 34788 5530 34790
rect 5554 34788 5610 34790
rect 5634 34788 5690 34790
rect 5394 33754 5450 33756
rect 5474 33754 5530 33756
rect 5554 33754 5610 33756
rect 5634 33754 5690 33756
rect 5394 33702 5440 33754
rect 5440 33702 5450 33754
rect 5474 33702 5504 33754
rect 5504 33702 5516 33754
rect 5516 33702 5530 33754
rect 5554 33702 5568 33754
rect 5568 33702 5580 33754
rect 5580 33702 5610 33754
rect 5634 33702 5644 33754
rect 5644 33702 5690 33754
rect 5394 33700 5450 33702
rect 5474 33700 5530 33702
rect 5554 33700 5610 33702
rect 5634 33700 5690 33702
rect 5394 32666 5450 32668
rect 5474 32666 5530 32668
rect 5554 32666 5610 32668
rect 5634 32666 5690 32668
rect 5394 32614 5440 32666
rect 5440 32614 5450 32666
rect 5474 32614 5504 32666
rect 5504 32614 5516 32666
rect 5516 32614 5530 32666
rect 5554 32614 5568 32666
rect 5568 32614 5580 32666
rect 5580 32614 5610 32666
rect 5634 32614 5644 32666
rect 5644 32614 5690 32666
rect 5394 32612 5450 32614
rect 5474 32612 5530 32614
rect 5554 32612 5610 32614
rect 5634 32612 5690 32614
rect 5394 31578 5450 31580
rect 5474 31578 5530 31580
rect 5554 31578 5610 31580
rect 5634 31578 5690 31580
rect 5394 31526 5440 31578
rect 5440 31526 5450 31578
rect 5474 31526 5504 31578
rect 5504 31526 5516 31578
rect 5516 31526 5530 31578
rect 5554 31526 5568 31578
rect 5568 31526 5580 31578
rect 5580 31526 5610 31578
rect 5634 31526 5644 31578
rect 5644 31526 5690 31578
rect 5394 31524 5450 31526
rect 5474 31524 5530 31526
rect 5554 31524 5610 31526
rect 5634 31524 5690 31526
rect 5394 30490 5450 30492
rect 5474 30490 5530 30492
rect 5554 30490 5610 30492
rect 5634 30490 5690 30492
rect 5394 30438 5440 30490
rect 5440 30438 5450 30490
rect 5474 30438 5504 30490
rect 5504 30438 5516 30490
rect 5516 30438 5530 30490
rect 5554 30438 5568 30490
rect 5568 30438 5580 30490
rect 5580 30438 5610 30490
rect 5634 30438 5644 30490
rect 5644 30438 5690 30490
rect 5394 30436 5450 30438
rect 5474 30436 5530 30438
rect 5554 30436 5610 30438
rect 5634 30436 5690 30438
rect 4710 30368 4766 30424
rect 3175 29946 3231 29948
rect 3255 29946 3311 29948
rect 3335 29946 3391 29948
rect 3415 29946 3471 29948
rect 3175 29894 3221 29946
rect 3221 29894 3231 29946
rect 3255 29894 3285 29946
rect 3285 29894 3297 29946
rect 3297 29894 3311 29946
rect 3335 29894 3349 29946
rect 3349 29894 3361 29946
rect 3361 29894 3391 29946
rect 3415 29894 3425 29946
rect 3425 29894 3471 29946
rect 3175 29892 3231 29894
rect 3255 29892 3311 29894
rect 3335 29892 3391 29894
rect 3415 29892 3471 29894
rect 3175 28858 3231 28860
rect 3255 28858 3311 28860
rect 3335 28858 3391 28860
rect 3415 28858 3471 28860
rect 3175 28806 3221 28858
rect 3221 28806 3231 28858
rect 3255 28806 3285 28858
rect 3285 28806 3297 28858
rect 3297 28806 3311 28858
rect 3335 28806 3349 28858
rect 3349 28806 3361 28858
rect 3361 28806 3391 28858
rect 3415 28806 3425 28858
rect 3425 28806 3471 28858
rect 3175 28804 3231 28806
rect 3255 28804 3311 28806
rect 3335 28804 3391 28806
rect 3415 28804 3471 28806
rect 3175 27770 3231 27772
rect 3255 27770 3311 27772
rect 3335 27770 3391 27772
rect 3415 27770 3471 27772
rect 3175 27718 3221 27770
rect 3221 27718 3231 27770
rect 3255 27718 3285 27770
rect 3285 27718 3297 27770
rect 3297 27718 3311 27770
rect 3335 27718 3349 27770
rect 3349 27718 3361 27770
rect 3361 27718 3391 27770
rect 3415 27718 3425 27770
rect 3425 27718 3471 27770
rect 3175 27716 3231 27718
rect 3255 27716 3311 27718
rect 3335 27716 3391 27718
rect 3415 27716 3471 27718
rect 2042 19352 2044 19372
rect 2044 19352 2096 19372
rect 2096 19352 2098 19372
rect 3175 26682 3231 26684
rect 3255 26682 3311 26684
rect 3335 26682 3391 26684
rect 3415 26682 3471 26684
rect 3175 26630 3221 26682
rect 3221 26630 3231 26682
rect 3255 26630 3285 26682
rect 3285 26630 3297 26682
rect 3297 26630 3311 26682
rect 3335 26630 3349 26682
rect 3349 26630 3361 26682
rect 3361 26630 3391 26682
rect 3415 26630 3425 26682
rect 3425 26630 3471 26682
rect 3175 26628 3231 26630
rect 3255 26628 3311 26630
rect 3335 26628 3391 26630
rect 3415 26628 3471 26630
rect 3175 25594 3231 25596
rect 3255 25594 3311 25596
rect 3335 25594 3391 25596
rect 3415 25594 3471 25596
rect 3175 25542 3221 25594
rect 3221 25542 3231 25594
rect 3255 25542 3285 25594
rect 3285 25542 3297 25594
rect 3297 25542 3311 25594
rect 3335 25542 3349 25594
rect 3349 25542 3361 25594
rect 3361 25542 3391 25594
rect 3415 25542 3425 25594
rect 3425 25542 3471 25594
rect 3175 25540 3231 25542
rect 3255 25540 3311 25542
rect 3335 25540 3391 25542
rect 3415 25540 3471 25542
rect 3175 24506 3231 24508
rect 3255 24506 3311 24508
rect 3335 24506 3391 24508
rect 3415 24506 3471 24508
rect 3175 24454 3221 24506
rect 3221 24454 3231 24506
rect 3255 24454 3285 24506
rect 3285 24454 3297 24506
rect 3297 24454 3311 24506
rect 3335 24454 3349 24506
rect 3349 24454 3361 24506
rect 3361 24454 3391 24506
rect 3415 24454 3425 24506
rect 3425 24454 3471 24506
rect 3175 24452 3231 24454
rect 3255 24452 3311 24454
rect 3335 24452 3391 24454
rect 3415 24452 3471 24454
rect 3175 23418 3231 23420
rect 3255 23418 3311 23420
rect 3335 23418 3391 23420
rect 3415 23418 3471 23420
rect 3175 23366 3221 23418
rect 3221 23366 3231 23418
rect 3255 23366 3285 23418
rect 3285 23366 3297 23418
rect 3297 23366 3311 23418
rect 3335 23366 3349 23418
rect 3349 23366 3361 23418
rect 3361 23366 3391 23418
rect 3415 23366 3425 23418
rect 3425 23366 3471 23418
rect 3175 23364 3231 23366
rect 3255 23364 3311 23366
rect 3335 23364 3391 23366
rect 3415 23364 3471 23366
rect 3175 22330 3231 22332
rect 3255 22330 3311 22332
rect 3335 22330 3391 22332
rect 3415 22330 3471 22332
rect 3175 22278 3221 22330
rect 3221 22278 3231 22330
rect 3255 22278 3285 22330
rect 3285 22278 3297 22330
rect 3297 22278 3311 22330
rect 3335 22278 3349 22330
rect 3349 22278 3361 22330
rect 3361 22278 3391 22330
rect 3415 22278 3425 22330
rect 3425 22278 3471 22330
rect 3175 22276 3231 22278
rect 3255 22276 3311 22278
rect 3335 22276 3391 22278
rect 3415 22276 3471 22278
rect 3175 21242 3231 21244
rect 3255 21242 3311 21244
rect 3335 21242 3391 21244
rect 3415 21242 3471 21244
rect 3175 21190 3221 21242
rect 3221 21190 3231 21242
rect 3255 21190 3285 21242
rect 3285 21190 3297 21242
rect 3297 21190 3311 21242
rect 3335 21190 3349 21242
rect 3349 21190 3361 21242
rect 3361 21190 3391 21242
rect 3415 21190 3425 21242
rect 3425 21190 3471 21242
rect 3175 21188 3231 21190
rect 3255 21188 3311 21190
rect 3335 21188 3391 21190
rect 3415 21188 3471 21190
rect 3175 20154 3231 20156
rect 3255 20154 3311 20156
rect 3335 20154 3391 20156
rect 3415 20154 3471 20156
rect 3175 20102 3221 20154
rect 3221 20102 3231 20154
rect 3255 20102 3285 20154
rect 3285 20102 3297 20154
rect 3297 20102 3311 20154
rect 3335 20102 3349 20154
rect 3349 20102 3361 20154
rect 3361 20102 3391 20154
rect 3415 20102 3425 20154
rect 3425 20102 3471 20154
rect 3175 20100 3231 20102
rect 3255 20100 3311 20102
rect 3335 20100 3391 20102
rect 3415 20100 3471 20102
rect 3175 19066 3231 19068
rect 3255 19066 3311 19068
rect 3335 19066 3391 19068
rect 3415 19066 3471 19068
rect 3175 19014 3221 19066
rect 3221 19014 3231 19066
rect 3255 19014 3285 19066
rect 3285 19014 3297 19066
rect 3297 19014 3311 19066
rect 3335 19014 3349 19066
rect 3349 19014 3361 19066
rect 3361 19014 3391 19066
rect 3415 19014 3425 19066
rect 3425 19014 3471 19066
rect 3175 19012 3231 19014
rect 3255 19012 3311 19014
rect 3335 19012 3391 19014
rect 3415 19012 3471 19014
rect 4250 27648 4306 27704
rect 5394 29402 5450 29404
rect 5474 29402 5530 29404
rect 5554 29402 5610 29404
rect 5634 29402 5690 29404
rect 5394 29350 5440 29402
rect 5440 29350 5450 29402
rect 5474 29350 5504 29402
rect 5504 29350 5516 29402
rect 5516 29350 5530 29402
rect 5554 29350 5568 29402
rect 5568 29350 5580 29402
rect 5580 29350 5610 29402
rect 5634 29350 5644 29402
rect 5644 29350 5690 29402
rect 5394 29348 5450 29350
rect 5474 29348 5530 29350
rect 5554 29348 5610 29350
rect 5634 29348 5690 29350
rect 4066 23432 4122 23488
rect 2778 12688 2834 12744
rect 2778 9696 2834 9752
rect 2686 6704 2742 6760
rect 2594 6432 2650 6488
rect 3175 17978 3231 17980
rect 3255 17978 3311 17980
rect 3335 17978 3391 17980
rect 3415 17978 3471 17980
rect 3175 17926 3221 17978
rect 3221 17926 3231 17978
rect 3255 17926 3285 17978
rect 3285 17926 3297 17978
rect 3297 17926 3311 17978
rect 3335 17926 3349 17978
rect 3349 17926 3361 17978
rect 3361 17926 3391 17978
rect 3415 17926 3425 17978
rect 3425 17926 3471 17978
rect 3175 17924 3231 17926
rect 3255 17924 3311 17926
rect 3335 17924 3391 17926
rect 3415 17924 3471 17926
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 3146 16652 3202 16688
rect 3146 16632 3148 16652
rect 3148 16632 3200 16652
rect 3200 16632 3202 16652
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 3606 12824 3662 12880
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 3606 11620 3662 11656
rect 3606 11600 3608 11620
rect 3608 11600 3660 11620
rect 3660 11600 3662 11620
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 3974 17196 4030 17232
rect 3974 17176 3976 17196
rect 3976 17176 4028 17196
rect 4028 17176 4030 17196
rect 4250 10920 4306 10976
rect 4066 9560 4122 9616
rect 5394 28314 5450 28316
rect 5474 28314 5530 28316
rect 5554 28314 5610 28316
rect 5634 28314 5690 28316
rect 5394 28262 5440 28314
rect 5440 28262 5450 28314
rect 5474 28262 5504 28314
rect 5504 28262 5516 28314
rect 5516 28262 5530 28314
rect 5554 28262 5568 28314
rect 5568 28262 5580 28314
rect 5580 28262 5610 28314
rect 5634 28262 5644 28314
rect 5644 28262 5690 28314
rect 5394 28260 5450 28262
rect 5474 28260 5530 28262
rect 5554 28260 5610 28262
rect 5634 28260 5690 28262
rect 5394 27226 5450 27228
rect 5474 27226 5530 27228
rect 5554 27226 5610 27228
rect 5634 27226 5690 27228
rect 5394 27174 5440 27226
rect 5440 27174 5450 27226
rect 5474 27174 5504 27226
rect 5504 27174 5516 27226
rect 5516 27174 5530 27226
rect 5554 27174 5568 27226
rect 5568 27174 5580 27226
rect 5580 27174 5610 27226
rect 5634 27174 5644 27226
rect 5644 27174 5690 27226
rect 5394 27172 5450 27174
rect 5474 27172 5530 27174
rect 5554 27172 5610 27174
rect 5634 27172 5690 27174
rect 5394 26138 5450 26140
rect 5474 26138 5530 26140
rect 5554 26138 5610 26140
rect 5634 26138 5690 26140
rect 5394 26086 5440 26138
rect 5440 26086 5450 26138
rect 5474 26086 5504 26138
rect 5504 26086 5516 26138
rect 5516 26086 5530 26138
rect 5554 26086 5568 26138
rect 5568 26086 5580 26138
rect 5580 26086 5610 26138
rect 5634 26086 5644 26138
rect 5644 26086 5690 26138
rect 5394 26084 5450 26086
rect 5474 26084 5530 26086
rect 5554 26084 5610 26086
rect 5634 26084 5690 26086
rect 5394 25050 5450 25052
rect 5474 25050 5530 25052
rect 5554 25050 5610 25052
rect 5634 25050 5690 25052
rect 5394 24998 5440 25050
rect 5440 24998 5450 25050
rect 5474 24998 5504 25050
rect 5504 24998 5516 25050
rect 5516 24998 5530 25050
rect 5554 24998 5568 25050
rect 5568 24998 5580 25050
rect 5580 24998 5610 25050
rect 5634 24998 5644 25050
rect 5644 24998 5690 25050
rect 5394 24996 5450 24998
rect 5474 24996 5530 24998
rect 5554 24996 5610 24998
rect 5634 24996 5690 24998
rect 5394 23962 5450 23964
rect 5474 23962 5530 23964
rect 5554 23962 5610 23964
rect 5634 23962 5690 23964
rect 5394 23910 5440 23962
rect 5440 23910 5450 23962
rect 5474 23910 5504 23962
rect 5504 23910 5516 23962
rect 5516 23910 5530 23962
rect 5554 23910 5568 23962
rect 5568 23910 5580 23962
rect 5580 23910 5610 23962
rect 5634 23910 5644 23962
rect 5644 23910 5690 23962
rect 5394 23908 5450 23910
rect 5474 23908 5530 23910
rect 5554 23908 5610 23910
rect 5634 23908 5690 23910
rect 5394 22874 5450 22876
rect 5474 22874 5530 22876
rect 5554 22874 5610 22876
rect 5634 22874 5690 22876
rect 5394 22822 5440 22874
rect 5440 22822 5450 22874
rect 5474 22822 5504 22874
rect 5504 22822 5516 22874
rect 5516 22822 5530 22874
rect 5554 22822 5568 22874
rect 5568 22822 5580 22874
rect 5580 22822 5610 22874
rect 5634 22822 5644 22874
rect 5644 22822 5690 22874
rect 5394 22820 5450 22822
rect 5474 22820 5530 22822
rect 5554 22820 5610 22822
rect 5634 22820 5690 22822
rect 9833 35930 9889 35932
rect 9913 35930 9969 35932
rect 9993 35930 10049 35932
rect 10073 35930 10129 35932
rect 9833 35878 9879 35930
rect 9879 35878 9889 35930
rect 9913 35878 9943 35930
rect 9943 35878 9955 35930
rect 9955 35878 9969 35930
rect 9993 35878 10007 35930
rect 10007 35878 10019 35930
rect 10019 35878 10049 35930
rect 10073 35878 10083 35930
rect 10083 35878 10129 35930
rect 9833 35876 9889 35878
rect 9913 35876 9969 35878
rect 9993 35876 10049 35878
rect 10073 35876 10129 35878
rect 14272 35930 14328 35932
rect 14352 35930 14408 35932
rect 14432 35930 14488 35932
rect 14512 35930 14568 35932
rect 14272 35878 14318 35930
rect 14318 35878 14328 35930
rect 14352 35878 14382 35930
rect 14382 35878 14394 35930
rect 14394 35878 14408 35930
rect 14432 35878 14446 35930
rect 14446 35878 14458 35930
rect 14458 35878 14488 35930
rect 14512 35878 14522 35930
rect 14522 35878 14568 35930
rect 14272 35876 14328 35878
rect 14352 35876 14408 35878
rect 14432 35876 14488 35878
rect 14512 35876 14568 35878
rect 18711 35930 18767 35932
rect 18791 35930 18847 35932
rect 18871 35930 18927 35932
rect 18951 35930 19007 35932
rect 18711 35878 18757 35930
rect 18757 35878 18767 35930
rect 18791 35878 18821 35930
rect 18821 35878 18833 35930
rect 18833 35878 18847 35930
rect 18871 35878 18885 35930
rect 18885 35878 18897 35930
rect 18897 35878 18927 35930
rect 18951 35878 18961 35930
rect 18961 35878 19007 35930
rect 18711 35876 18767 35878
rect 18791 35876 18847 35878
rect 18871 35876 18927 35878
rect 18951 35876 19007 35878
rect 7614 35386 7670 35388
rect 7694 35386 7750 35388
rect 7774 35386 7830 35388
rect 7854 35386 7910 35388
rect 7614 35334 7660 35386
rect 7660 35334 7670 35386
rect 7694 35334 7724 35386
rect 7724 35334 7736 35386
rect 7736 35334 7750 35386
rect 7774 35334 7788 35386
rect 7788 35334 7800 35386
rect 7800 35334 7830 35386
rect 7854 35334 7864 35386
rect 7864 35334 7910 35386
rect 7614 35332 7670 35334
rect 7694 35332 7750 35334
rect 7774 35332 7830 35334
rect 7854 35332 7910 35334
rect 12053 35386 12109 35388
rect 12133 35386 12189 35388
rect 12213 35386 12269 35388
rect 12293 35386 12349 35388
rect 12053 35334 12099 35386
rect 12099 35334 12109 35386
rect 12133 35334 12163 35386
rect 12163 35334 12175 35386
rect 12175 35334 12189 35386
rect 12213 35334 12227 35386
rect 12227 35334 12239 35386
rect 12239 35334 12269 35386
rect 12293 35334 12303 35386
rect 12303 35334 12349 35386
rect 12053 35332 12109 35334
rect 12133 35332 12189 35334
rect 12213 35332 12269 35334
rect 12293 35332 12349 35334
rect 16492 35386 16548 35388
rect 16572 35386 16628 35388
rect 16652 35386 16708 35388
rect 16732 35386 16788 35388
rect 16492 35334 16538 35386
rect 16538 35334 16548 35386
rect 16572 35334 16602 35386
rect 16602 35334 16614 35386
rect 16614 35334 16628 35386
rect 16652 35334 16666 35386
rect 16666 35334 16678 35386
rect 16678 35334 16708 35386
rect 16732 35334 16742 35386
rect 16742 35334 16788 35386
rect 16492 35332 16548 35334
rect 16572 35332 16628 35334
rect 16652 35332 16708 35334
rect 16732 35332 16788 35334
rect 9833 34842 9889 34844
rect 9913 34842 9969 34844
rect 9993 34842 10049 34844
rect 10073 34842 10129 34844
rect 9833 34790 9879 34842
rect 9879 34790 9889 34842
rect 9913 34790 9943 34842
rect 9943 34790 9955 34842
rect 9955 34790 9969 34842
rect 9993 34790 10007 34842
rect 10007 34790 10019 34842
rect 10019 34790 10049 34842
rect 10073 34790 10083 34842
rect 10083 34790 10129 34842
rect 9833 34788 9889 34790
rect 9913 34788 9969 34790
rect 9993 34788 10049 34790
rect 10073 34788 10129 34790
rect 14272 34842 14328 34844
rect 14352 34842 14408 34844
rect 14432 34842 14488 34844
rect 14512 34842 14568 34844
rect 14272 34790 14318 34842
rect 14318 34790 14328 34842
rect 14352 34790 14382 34842
rect 14382 34790 14394 34842
rect 14394 34790 14408 34842
rect 14432 34790 14446 34842
rect 14446 34790 14458 34842
rect 14458 34790 14488 34842
rect 14512 34790 14522 34842
rect 14522 34790 14568 34842
rect 14272 34788 14328 34790
rect 14352 34788 14408 34790
rect 14432 34788 14488 34790
rect 14512 34788 14568 34790
rect 18711 34842 18767 34844
rect 18791 34842 18847 34844
rect 18871 34842 18927 34844
rect 18951 34842 19007 34844
rect 18711 34790 18757 34842
rect 18757 34790 18767 34842
rect 18791 34790 18821 34842
rect 18821 34790 18833 34842
rect 18833 34790 18847 34842
rect 18871 34790 18885 34842
rect 18885 34790 18897 34842
rect 18897 34790 18927 34842
rect 18951 34790 18961 34842
rect 18961 34790 19007 34842
rect 18711 34788 18767 34790
rect 18791 34788 18847 34790
rect 18871 34788 18927 34790
rect 18951 34788 19007 34790
rect 7614 34298 7670 34300
rect 7694 34298 7750 34300
rect 7774 34298 7830 34300
rect 7854 34298 7910 34300
rect 7614 34246 7660 34298
rect 7660 34246 7670 34298
rect 7694 34246 7724 34298
rect 7724 34246 7736 34298
rect 7736 34246 7750 34298
rect 7774 34246 7788 34298
rect 7788 34246 7800 34298
rect 7800 34246 7830 34298
rect 7854 34246 7864 34298
rect 7864 34246 7910 34298
rect 7614 34244 7670 34246
rect 7694 34244 7750 34246
rect 7774 34244 7830 34246
rect 7854 34244 7910 34246
rect 12053 34298 12109 34300
rect 12133 34298 12189 34300
rect 12213 34298 12269 34300
rect 12293 34298 12349 34300
rect 12053 34246 12099 34298
rect 12099 34246 12109 34298
rect 12133 34246 12163 34298
rect 12163 34246 12175 34298
rect 12175 34246 12189 34298
rect 12213 34246 12227 34298
rect 12227 34246 12239 34298
rect 12239 34246 12269 34298
rect 12293 34246 12303 34298
rect 12303 34246 12349 34298
rect 12053 34244 12109 34246
rect 12133 34244 12189 34246
rect 12213 34244 12269 34246
rect 12293 34244 12349 34246
rect 16492 34298 16548 34300
rect 16572 34298 16628 34300
rect 16652 34298 16708 34300
rect 16732 34298 16788 34300
rect 16492 34246 16538 34298
rect 16538 34246 16548 34298
rect 16572 34246 16602 34298
rect 16602 34246 16614 34298
rect 16614 34246 16628 34298
rect 16652 34246 16666 34298
rect 16666 34246 16678 34298
rect 16678 34246 16708 34298
rect 16732 34246 16742 34298
rect 16742 34246 16788 34298
rect 16492 34244 16548 34246
rect 16572 34244 16628 34246
rect 16652 34244 16708 34246
rect 16732 34244 16788 34246
rect 5394 21786 5450 21788
rect 5474 21786 5530 21788
rect 5554 21786 5610 21788
rect 5634 21786 5690 21788
rect 5394 21734 5440 21786
rect 5440 21734 5450 21786
rect 5474 21734 5504 21786
rect 5504 21734 5516 21786
rect 5516 21734 5530 21786
rect 5554 21734 5568 21786
rect 5568 21734 5580 21786
rect 5580 21734 5610 21786
rect 5634 21734 5644 21786
rect 5644 21734 5690 21786
rect 5394 21732 5450 21734
rect 5474 21732 5530 21734
rect 5554 21732 5610 21734
rect 5634 21732 5690 21734
rect 6182 26308 6238 26344
rect 6182 26288 6184 26308
rect 6184 26288 6236 26308
rect 6236 26288 6238 26308
rect 5394 20698 5450 20700
rect 5474 20698 5530 20700
rect 5554 20698 5610 20700
rect 5634 20698 5690 20700
rect 5394 20646 5440 20698
rect 5440 20646 5450 20698
rect 5474 20646 5504 20698
rect 5504 20646 5516 20698
rect 5516 20646 5530 20698
rect 5554 20646 5568 20698
rect 5568 20646 5580 20698
rect 5580 20646 5610 20698
rect 5634 20646 5644 20698
rect 5644 20646 5690 20698
rect 5394 20644 5450 20646
rect 5474 20644 5530 20646
rect 5554 20644 5610 20646
rect 5634 20644 5690 20646
rect 4802 5480 4858 5536
rect 5394 19610 5450 19612
rect 5474 19610 5530 19612
rect 5554 19610 5610 19612
rect 5634 19610 5690 19612
rect 5394 19558 5440 19610
rect 5440 19558 5450 19610
rect 5474 19558 5504 19610
rect 5504 19558 5516 19610
rect 5516 19558 5530 19610
rect 5554 19558 5568 19610
rect 5568 19558 5580 19610
rect 5580 19558 5610 19610
rect 5634 19558 5644 19610
rect 5644 19558 5690 19610
rect 5394 19556 5450 19558
rect 5474 19556 5530 19558
rect 5554 19556 5610 19558
rect 5634 19556 5690 19558
rect 5394 18522 5450 18524
rect 5474 18522 5530 18524
rect 5554 18522 5610 18524
rect 5634 18522 5690 18524
rect 5394 18470 5440 18522
rect 5440 18470 5450 18522
rect 5474 18470 5504 18522
rect 5504 18470 5516 18522
rect 5516 18470 5530 18522
rect 5554 18470 5568 18522
rect 5568 18470 5580 18522
rect 5580 18470 5610 18522
rect 5634 18470 5644 18522
rect 5644 18470 5690 18522
rect 5394 18468 5450 18470
rect 5474 18468 5530 18470
rect 5554 18468 5610 18470
rect 5634 18468 5690 18470
rect 5394 17434 5450 17436
rect 5474 17434 5530 17436
rect 5554 17434 5610 17436
rect 5634 17434 5690 17436
rect 5394 17382 5440 17434
rect 5440 17382 5450 17434
rect 5474 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5530 17434
rect 5554 17382 5568 17434
rect 5568 17382 5580 17434
rect 5580 17382 5610 17434
rect 5634 17382 5644 17434
rect 5644 17382 5690 17434
rect 5394 17380 5450 17382
rect 5474 17380 5530 17382
rect 5554 17380 5610 17382
rect 5634 17380 5690 17382
rect 5394 16346 5450 16348
rect 5474 16346 5530 16348
rect 5554 16346 5610 16348
rect 5634 16346 5690 16348
rect 5394 16294 5440 16346
rect 5440 16294 5450 16346
rect 5474 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5530 16346
rect 5554 16294 5568 16346
rect 5568 16294 5580 16346
rect 5580 16294 5610 16346
rect 5634 16294 5644 16346
rect 5644 16294 5690 16346
rect 5394 16292 5450 16294
rect 5474 16292 5530 16294
rect 5554 16292 5610 16294
rect 5634 16292 5690 16294
rect 938 1944 994 2000
rect 5394 15258 5450 15260
rect 5474 15258 5530 15260
rect 5554 15258 5610 15260
rect 5634 15258 5690 15260
rect 5394 15206 5440 15258
rect 5440 15206 5450 15258
rect 5474 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5530 15258
rect 5554 15206 5568 15258
rect 5568 15206 5580 15258
rect 5580 15206 5610 15258
rect 5634 15206 5644 15258
rect 5644 15206 5690 15258
rect 5394 15204 5450 15206
rect 5474 15204 5530 15206
rect 5554 15204 5610 15206
rect 5634 15204 5690 15206
rect 5394 14170 5450 14172
rect 5474 14170 5530 14172
rect 5554 14170 5610 14172
rect 5634 14170 5690 14172
rect 5394 14118 5440 14170
rect 5440 14118 5450 14170
rect 5474 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5530 14170
rect 5554 14118 5568 14170
rect 5568 14118 5580 14170
rect 5580 14118 5610 14170
rect 5634 14118 5644 14170
rect 5644 14118 5690 14170
rect 5394 14116 5450 14118
rect 5474 14116 5530 14118
rect 5554 14116 5610 14118
rect 5634 14116 5690 14118
rect 5170 13776 5226 13832
rect 5394 13082 5450 13084
rect 5474 13082 5530 13084
rect 5554 13082 5610 13084
rect 5634 13082 5690 13084
rect 5394 13030 5440 13082
rect 5440 13030 5450 13082
rect 5474 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5530 13082
rect 5554 13030 5568 13082
rect 5568 13030 5580 13082
rect 5580 13030 5610 13082
rect 5634 13030 5644 13082
rect 5644 13030 5690 13082
rect 5394 13028 5450 13030
rect 5474 13028 5530 13030
rect 5554 13028 5610 13030
rect 5634 13028 5690 13030
rect 5394 11994 5450 11996
rect 5474 11994 5530 11996
rect 5554 11994 5610 11996
rect 5634 11994 5690 11996
rect 5394 11942 5440 11994
rect 5440 11942 5450 11994
rect 5474 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5530 11994
rect 5554 11942 5568 11994
rect 5568 11942 5580 11994
rect 5580 11942 5610 11994
rect 5634 11942 5644 11994
rect 5644 11942 5690 11994
rect 5394 11940 5450 11942
rect 5474 11940 5530 11942
rect 5554 11940 5610 11942
rect 5634 11940 5690 11942
rect 5394 10906 5450 10908
rect 5474 10906 5530 10908
rect 5554 10906 5610 10908
rect 5634 10906 5690 10908
rect 5394 10854 5440 10906
rect 5440 10854 5450 10906
rect 5474 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5530 10906
rect 5554 10854 5568 10906
rect 5568 10854 5580 10906
rect 5580 10854 5610 10906
rect 5634 10854 5644 10906
rect 5644 10854 5690 10906
rect 5394 10852 5450 10854
rect 5474 10852 5530 10854
rect 5554 10852 5610 10854
rect 5634 10852 5690 10854
rect 5394 9818 5450 9820
rect 5474 9818 5530 9820
rect 5554 9818 5610 9820
rect 5634 9818 5690 9820
rect 5394 9766 5440 9818
rect 5440 9766 5450 9818
rect 5474 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5530 9818
rect 5554 9766 5568 9818
rect 5568 9766 5580 9818
rect 5580 9766 5610 9818
rect 5634 9766 5644 9818
rect 5644 9766 5690 9818
rect 5394 9764 5450 9766
rect 5474 9764 5530 9766
rect 5554 9764 5610 9766
rect 5634 9764 5690 9766
rect 5394 8730 5450 8732
rect 5474 8730 5530 8732
rect 5554 8730 5610 8732
rect 5634 8730 5690 8732
rect 5394 8678 5440 8730
rect 5440 8678 5450 8730
rect 5474 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5530 8730
rect 5554 8678 5568 8730
rect 5568 8678 5580 8730
rect 5580 8678 5610 8730
rect 5634 8678 5644 8730
rect 5644 8678 5690 8730
rect 5394 8676 5450 8678
rect 5474 8676 5530 8678
rect 5554 8676 5610 8678
rect 5634 8676 5690 8678
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 6826 20712 6882 20768
rect 7010 24112 7066 24168
rect 6826 6568 6882 6624
rect 7614 33210 7670 33212
rect 7694 33210 7750 33212
rect 7774 33210 7830 33212
rect 7854 33210 7910 33212
rect 7614 33158 7660 33210
rect 7660 33158 7670 33210
rect 7694 33158 7724 33210
rect 7724 33158 7736 33210
rect 7736 33158 7750 33210
rect 7774 33158 7788 33210
rect 7788 33158 7800 33210
rect 7800 33158 7830 33210
rect 7854 33158 7864 33210
rect 7864 33158 7910 33210
rect 7614 33156 7670 33158
rect 7694 33156 7750 33158
rect 7774 33156 7830 33158
rect 7854 33156 7910 33158
rect 7614 32122 7670 32124
rect 7694 32122 7750 32124
rect 7774 32122 7830 32124
rect 7854 32122 7910 32124
rect 7614 32070 7660 32122
rect 7660 32070 7670 32122
rect 7694 32070 7724 32122
rect 7724 32070 7736 32122
rect 7736 32070 7750 32122
rect 7774 32070 7788 32122
rect 7788 32070 7800 32122
rect 7800 32070 7830 32122
rect 7854 32070 7864 32122
rect 7864 32070 7910 32122
rect 7614 32068 7670 32070
rect 7694 32068 7750 32070
rect 7774 32068 7830 32070
rect 7854 32068 7910 32070
rect 7614 31034 7670 31036
rect 7694 31034 7750 31036
rect 7774 31034 7830 31036
rect 7854 31034 7910 31036
rect 7614 30982 7660 31034
rect 7660 30982 7670 31034
rect 7694 30982 7724 31034
rect 7724 30982 7736 31034
rect 7736 30982 7750 31034
rect 7774 30982 7788 31034
rect 7788 30982 7800 31034
rect 7800 30982 7830 31034
rect 7854 30982 7864 31034
rect 7864 30982 7910 31034
rect 7614 30980 7670 30982
rect 7694 30980 7750 30982
rect 7774 30980 7830 30982
rect 7854 30980 7910 30982
rect 7614 29946 7670 29948
rect 7694 29946 7750 29948
rect 7774 29946 7830 29948
rect 7854 29946 7910 29948
rect 7614 29894 7660 29946
rect 7660 29894 7670 29946
rect 7694 29894 7724 29946
rect 7724 29894 7736 29946
rect 7736 29894 7750 29946
rect 7774 29894 7788 29946
rect 7788 29894 7800 29946
rect 7800 29894 7830 29946
rect 7854 29894 7864 29946
rect 7864 29894 7910 29946
rect 7614 29892 7670 29894
rect 7694 29892 7750 29894
rect 7774 29892 7830 29894
rect 7854 29892 7910 29894
rect 7614 28858 7670 28860
rect 7694 28858 7750 28860
rect 7774 28858 7830 28860
rect 7854 28858 7910 28860
rect 7614 28806 7660 28858
rect 7660 28806 7670 28858
rect 7694 28806 7724 28858
rect 7724 28806 7736 28858
rect 7736 28806 7750 28858
rect 7774 28806 7788 28858
rect 7788 28806 7800 28858
rect 7800 28806 7830 28858
rect 7854 28806 7864 28858
rect 7864 28806 7910 28858
rect 7614 28804 7670 28806
rect 7694 28804 7750 28806
rect 7774 28804 7830 28806
rect 7854 28804 7910 28806
rect 7614 27770 7670 27772
rect 7694 27770 7750 27772
rect 7774 27770 7830 27772
rect 7854 27770 7910 27772
rect 7614 27718 7660 27770
rect 7660 27718 7670 27770
rect 7694 27718 7724 27770
rect 7724 27718 7736 27770
rect 7736 27718 7750 27770
rect 7774 27718 7788 27770
rect 7788 27718 7800 27770
rect 7800 27718 7830 27770
rect 7854 27718 7864 27770
rect 7864 27718 7910 27770
rect 7614 27716 7670 27718
rect 7694 27716 7750 27718
rect 7774 27716 7830 27718
rect 7854 27716 7910 27718
rect 7470 27104 7526 27160
rect 7614 26682 7670 26684
rect 7694 26682 7750 26684
rect 7774 26682 7830 26684
rect 7854 26682 7910 26684
rect 7614 26630 7660 26682
rect 7660 26630 7670 26682
rect 7694 26630 7724 26682
rect 7724 26630 7736 26682
rect 7736 26630 7750 26682
rect 7774 26630 7788 26682
rect 7788 26630 7800 26682
rect 7800 26630 7830 26682
rect 7854 26630 7864 26682
rect 7864 26630 7910 26682
rect 7614 26628 7670 26630
rect 7694 26628 7750 26630
rect 7774 26628 7830 26630
rect 7854 26628 7910 26630
rect 8114 29008 8170 29064
rect 7614 25594 7670 25596
rect 7694 25594 7750 25596
rect 7774 25594 7830 25596
rect 7854 25594 7910 25596
rect 7614 25542 7660 25594
rect 7660 25542 7670 25594
rect 7694 25542 7724 25594
rect 7724 25542 7736 25594
rect 7736 25542 7750 25594
rect 7774 25542 7788 25594
rect 7788 25542 7800 25594
rect 7800 25542 7830 25594
rect 7854 25542 7864 25594
rect 7864 25542 7910 25594
rect 7614 25540 7670 25542
rect 7694 25540 7750 25542
rect 7774 25540 7830 25542
rect 7854 25540 7910 25542
rect 7838 25236 7840 25256
rect 7840 25236 7892 25256
rect 7892 25236 7894 25256
rect 7838 25200 7894 25236
rect 7614 24506 7670 24508
rect 7694 24506 7750 24508
rect 7774 24506 7830 24508
rect 7854 24506 7910 24508
rect 7614 24454 7660 24506
rect 7660 24454 7670 24506
rect 7694 24454 7724 24506
rect 7724 24454 7736 24506
rect 7736 24454 7750 24506
rect 7774 24454 7788 24506
rect 7788 24454 7800 24506
rect 7800 24454 7830 24506
rect 7854 24454 7864 24506
rect 7864 24454 7910 24506
rect 7614 24452 7670 24454
rect 7694 24452 7750 24454
rect 7774 24452 7830 24454
rect 7854 24452 7910 24454
rect 7614 23418 7670 23420
rect 7694 23418 7750 23420
rect 7774 23418 7830 23420
rect 7854 23418 7910 23420
rect 7614 23366 7660 23418
rect 7660 23366 7670 23418
rect 7694 23366 7724 23418
rect 7724 23366 7736 23418
rect 7736 23366 7750 23418
rect 7774 23366 7788 23418
rect 7788 23366 7800 23418
rect 7800 23366 7830 23418
rect 7854 23366 7864 23418
rect 7864 23366 7910 23418
rect 7614 23364 7670 23366
rect 7694 23364 7750 23366
rect 7774 23364 7830 23366
rect 7854 23364 7910 23366
rect 7614 22330 7670 22332
rect 7694 22330 7750 22332
rect 7774 22330 7830 22332
rect 7854 22330 7910 22332
rect 7614 22278 7660 22330
rect 7660 22278 7670 22330
rect 7694 22278 7724 22330
rect 7724 22278 7736 22330
rect 7736 22278 7750 22330
rect 7774 22278 7788 22330
rect 7788 22278 7800 22330
rect 7800 22278 7830 22330
rect 7854 22278 7864 22330
rect 7864 22278 7910 22330
rect 7614 22276 7670 22278
rect 7694 22276 7750 22278
rect 7774 22276 7830 22278
rect 7854 22276 7910 22278
rect 7614 21242 7670 21244
rect 7694 21242 7750 21244
rect 7774 21242 7830 21244
rect 7854 21242 7910 21244
rect 7614 21190 7660 21242
rect 7660 21190 7670 21242
rect 7694 21190 7724 21242
rect 7724 21190 7736 21242
rect 7736 21190 7750 21242
rect 7774 21190 7788 21242
rect 7788 21190 7800 21242
rect 7800 21190 7830 21242
rect 7854 21190 7864 21242
rect 7864 21190 7910 21242
rect 7614 21188 7670 21190
rect 7694 21188 7750 21190
rect 7774 21188 7830 21190
rect 7854 21188 7910 21190
rect 7614 20154 7670 20156
rect 7694 20154 7750 20156
rect 7774 20154 7830 20156
rect 7854 20154 7910 20156
rect 7614 20102 7660 20154
rect 7660 20102 7670 20154
rect 7694 20102 7724 20154
rect 7724 20102 7736 20154
rect 7736 20102 7750 20154
rect 7774 20102 7788 20154
rect 7788 20102 7800 20154
rect 7800 20102 7830 20154
rect 7854 20102 7864 20154
rect 7864 20102 7910 20154
rect 7614 20100 7670 20102
rect 7694 20100 7750 20102
rect 7774 20100 7830 20102
rect 7854 20100 7910 20102
rect 7614 19066 7670 19068
rect 7694 19066 7750 19068
rect 7774 19066 7830 19068
rect 7854 19066 7910 19068
rect 7614 19014 7660 19066
rect 7660 19014 7670 19066
rect 7694 19014 7724 19066
rect 7724 19014 7736 19066
rect 7736 19014 7750 19066
rect 7774 19014 7788 19066
rect 7788 19014 7800 19066
rect 7800 19014 7830 19066
rect 7854 19014 7864 19066
rect 7864 19014 7910 19066
rect 7614 19012 7670 19014
rect 7694 19012 7750 19014
rect 7774 19012 7830 19014
rect 7854 19012 7910 19014
rect 7614 17978 7670 17980
rect 7694 17978 7750 17980
rect 7774 17978 7830 17980
rect 7854 17978 7910 17980
rect 7614 17926 7660 17978
rect 7660 17926 7670 17978
rect 7694 17926 7724 17978
rect 7724 17926 7736 17978
rect 7736 17926 7750 17978
rect 7774 17926 7788 17978
rect 7788 17926 7800 17978
rect 7800 17926 7830 17978
rect 7854 17926 7864 17978
rect 7864 17926 7910 17978
rect 7614 17924 7670 17926
rect 7694 17924 7750 17926
rect 7774 17924 7830 17926
rect 7854 17924 7910 17926
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 9833 33754 9889 33756
rect 9913 33754 9969 33756
rect 9993 33754 10049 33756
rect 10073 33754 10129 33756
rect 9833 33702 9879 33754
rect 9879 33702 9889 33754
rect 9913 33702 9943 33754
rect 9943 33702 9955 33754
rect 9955 33702 9969 33754
rect 9993 33702 10007 33754
rect 10007 33702 10019 33754
rect 10019 33702 10049 33754
rect 10073 33702 10083 33754
rect 10083 33702 10129 33754
rect 9833 33700 9889 33702
rect 9913 33700 9969 33702
rect 9993 33700 10049 33702
rect 10073 33700 10129 33702
rect 14272 33754 14328 33756
rect 14352 33754 14408 33756
rect 14432 33754 14488 33756
rect 14512 33754 14568 33756
rect 14272 33702 14318 33754
rect 14318 33702 14328 33754
rect 14352 33702 14382 33754
rect 14382 33702 14394 33754
rect 14394 33702 14408 33754
rect 14432 33702 14446 33754
rect 14446 33702 14458 33754
rect 14458 33702 14488 33754
rect 14512 33702 14522 33754
rect 14522 33702 14568 33754
rect 14272 33700 14328 33702
rect 14352 33700 14408 33702
rect 14432 33700 14488 33702
rect 14512 33700 14568 33702
rect 18711 33754 18767 33756
rect 18791 33754 18847 33756
rect 18871 33754 18927 33756
rect 18951 33754 19007 33756
rect 18711 33702 18757 33754
rect 18757 33702 18767 33754
rect 18791 33702 18821 33754
rect 18821 33702 18833 33754
rect 18833 33702 18847 33754
rect 18871 33702 18885 33754
rect 18885 33702 18897 33754
rect 18897 33702 18927 33754
rect 18951 33702 18961 33754
rect 18961 33702 19007 33754
rect 18711 33700 18767 33702
rect 18791 33700 18847 33702
rect 18871 33700 18927 33702
rect 18951 33700 19007 33702
rect 12053 33210 12109 33212
rect 12133 33210 12189 33212
rect 12213 33210 12269 33212
rect 12293 33210 12349 33212
rect 12053 33158 12099 33210
rect 12099 33158 12109 33210
rect 12133 33158 12163 33210
rect 12163 33158 12175 33210
rect 12175 33158 12189 33210
rect 12213 33158 12227 33210
rect 12227 33158 12239 33210
rect 12239 33158 12269 33210
rect 12293 33158 12303 33210
rect 12303 33158 12349 33210
rect 12053 33156 12109 33158
rect 12133 33156 12189 33158
rect 12213 33156 12269 33158
rect 12293 33156 12349 33158
rect 16492 33210 16548 33212
rect 16572 33210 16628 33212
rect 16652 33210 16708 33212
rect 16732 33210 16788 33212
rect 16492 33158 16538 33210
rect 16538 33158 16548 33210
rect 16572 33158 16602 33210
rect 16602 33158 16614 33210
rect 16614 33158 16628 33210
rect 16652 33158 16666 33210
rect 16666 33158 16678 33210
rect 16678 33158 16708 33210
rect 16732 33158 16742 33210
rect 16742 33158 16788 33210
rect 16492 33156 16548 33158
rect 16572 33156 16628 33158
rect 16652 33156 16708 33158
rect 16732 33156 16788 33158
rect 9833 32666 9889 32668
rect 9913 32666 9969 32668
rect 9993 32666 10049 32668
rect 10073 32666 10129 32668
rect 9833 32614 9879 32666
rect 9879 32614 9889 32666
rect 9913 32614 9943 32666
rect 9943 32614 9955 32666
rect 9955 32614 9969 32666
rect 9993 32614 10007 32666
rect 10007 32614 10019 32666
rect 10019 32614 10049 32666
rect 10073 32614 10083 32666
rect 10083 32614 10129 32666
rect 9833 32612 9889 32614
rect 9913 32612 9969 32614
rect 9993 32612 10049 32614
rect 10073 32612 10129 32614
rect 14272 32666 14328 32668
rect 14352 32666 14408 32668
rect 14432 32666 14488 32668
rect 14512 32666 14568 32668
rect 14272 32614 14318 32666
rect 14318 32614 14328 32666
rect 14352 32614 14382 32666
rect 14382 32614 14394 32666
rect 14394 32614 14408 32666
rect 14432 32614 14446 32666
rect 14446 32614 14458 32666
rect 14458 32614 14488 32666
rect 14512 32614 14522 32666
rect 14522 32614 14568 32666
rect 14272 32612 14328 32614
rect 14352 32612 14408 32614
rect 14432 32612 14488 32614
rect 14512 32612 14568 32614
rect 18711 32666 18767 32668
rect 18791 32666 18847 32668
rect 18871 32666 18927 32668
rect 18951 32666 19007 32668
rect 18711 32614 18757 32666
rect 18757 32614 18767 32666
rect 18791 32614 18821 32666
rect 18821 32614 18833 32666
rect 18833 32614 18847 32666
rect 18871 32614 18885 32666
rect 18885 32614 18897 32666
rect 18897 32614 18927 32666
rect 18951 32614 18961 32666
rect 18961 32614 19007 32666
rect 18711 32612 18767 32614
rect 18791 32612 18847 32614
rect 18871 32612 18927 32614
rect 18951 32612 19007 32614
rect 12053 32122 12109 32124
rect 12133 32122 12189 32124
rect 12213 32122 12269 32124
rect 12293 32122 12349 32124
rect 12053 32070 12099 32122
rect 12099 32070 12109 32122
rect 12133 32070 12163 32122
rect 12163 32070 12175 32122
rect 12175 32070 12189 32122
rect 12213 32070 12227 32122
rect 12227 32070 12239 32122
rect 12239 32070 12269 32122
rect 12293 32070 12303 32122
rect 12303 32070 12349 32122
rect 12053 32068 12109 32070
rect 12133 32068 12189 32070
rect 12213 32068 12269 32070
rect 12293 32068 12349 32070
rect 16492 32122 16548 32124
rect 16572 32122 16628 32124
rect 16652 32122 16708 32124
rect 16732 32122 16788 32124
rect 16492 32070 16538 32122
rect 16538 32070 16548 32122
rect 16572 32070 16602 32122
rect 16602 32070 16614 32122
rect 16614 32070 16628 32122
rect 16652 32070 16666 32122
rect 16666 32070 16678 32122
rect 16678 32070 16708 32122
rect 16732 32070 16742 32122
rect 16742 32070 16788 32122
rect 16492 32068 16548 32070
rect 16572 32068 16628 32070
rect 16652 32068 16708 32070
rect 16732 32068 16788 32070
rect 9833 31578 9889 31580
rect 9913 31578 9969 31580
rect 9993 31578 10049 31580
rect 10073 31578 10129 31580
rect 9833 31526 9879 31578
rect 9879 31526 9889 31578
rect 9913 31526 9943 31578
rect 9943 31526 9955 31578
rect 9955 31526 9969 31578
rect 9993 31526 10007 31578
rect 10007 31526 10019 31578
rect 10019 31526 10049 31578
rect 10073 31526 10083 31578
rect 10083 31526 10129 31578
rect 9833 31524 9889 31526
rect 9913 31524 9969 31526
rect 9993 31524 10049 31526
rect 10073 31524 10129 31526
rect 14272 31578 14328 31580
rect 14352 31578 14408 31580
rect 14432 31578 14488 31580
rect 14512 31578 14568 31580
rect 14272 31526 14318 31578
rect 14318 31526 14328 31578
rect 14352 31526 14382 31578
rect 14382 31526 14394 31578
rect 14394 31526 14408 31578
rect 14432 31526 14446 31578
rect 14446 31526 14458 31578
rect 14458 31526 14488 31578
rect 14512 31526 14522 31578
rect 14522 31526 14568 31578
rect 14272 31524 14328 31526
rect 14352 31524 14408 31526
rect 14432 31524 14488 31526
rect 14512 31524 14568 31526
rect 18711 31578 18767 31580
rect 18791 31578 18847 31580
rect 18871 31578 18927 31580
rect 18951 31578 19007 31580
rect 18711 31526 18757 31578
rect 18757 31526 18767 31578
rect 18791 31526 18821 31578
rect 18821 31526 18833 31578
rect 18833 31526 18847 31578
rect 18871 31526 18885 31578
rect 18885 31526 18897 31578
rect 18897 31526 18927 31578
rect 18951 31526 18961 31578
rect 18961 31526 19007 31578
rect 18711 31524 18767 31526
rect 18791 31524 18847 31526
rect 18871 31524 18927 31526
rect 18951 31524 19007 31526
rect 12053 31034 12109 31036
rect 12133 31034 12189 31036
rect 12213 31034 12269 31036
rect 12293 31034 12349 31036
rect 12053 30982 12099 31034
rect 12099 30982 12109 31034
rect 12133 30982 12163 31034
rect 12163 30982 12175 31034
rect 12175 30982 12189 31034
rect 12213 30982 12227 31034
rect 12227 30982 12239 31034
rect 12239 30982 12269 31034
rect 12293 30982 12303 31034
rect 12303 30982 12349 31034
rect 12053 30980 12109 30982
rect 12133 30980 12189 30982
rect 12213 30980 12269 30982
rect 12293 30980 12349 30982
rect 16492 31034 16548 31036
rect 16572 31034 16628 31036
rect 16652 31034 16708 31036
rect 16732 31034 16788 31036
rect 16492 30982 16538 31034
rect 16538 30982 16548 31034
rect 16572 30982 16602 31034
rect 16602 30982 16614 31034
rect 16614 30982 16628 31034
rect 16652 30982 16666 31034
rect 16666 30982 16678 31034
rect 16678 30982 16708 31034
rect 16732 30982 16742 31034
rect 16742 30982 16788 31034
rect 16492 30980 16548 30982
rect 16572 30980 16628 30982
rect 16652 30980 16708 30982
rect 16732 30980 16788 30982
rect 9833 30490 9889 30492
rect 9913 30490 9969 30492
rect 9993 30490 10049 30492
rect 10073 30490 10129 30492
rect 9833 30438 9879 30490
rect 9879 30438 9889 30490
rect 9913 30438 9943 30490
rect 9943 30438 9955 30490
rect 9955 30438 9969 30490
rect 9993 30438 10007 30490
rect 10007 30438 10019 30490
rect 10019 30438 10049 30490
rect 10073 30438 10083 30490
rect 10083 30438 10129 30490
rect 9833 30436 9889 30438
rect 9913 30436 9969 30438
rect 9993 30436 10049 30438
rect 10073 30436 10129 30438
rect 14272 30490 14328 30492
rect 14352 30490 14408 30492
rect 14432 30490 14488 30492
rect 14512 30490 14568 30492
rect 14272 30438 14318 30490
rect 14318 30438 14328 30490
rect 14352 30438 14382 30490
rect 14382 30438 14394 30490
rect 14394 30438 14408 30490
rect 14432 30438 14446 30490
rect 14446 30438 14458 30490
rect 14458 30438 14488 30490
rect 14512 30438 14522 30490
rect 14522 30438 14568 30490
rect 14272 30436 14328 30438
rect 14352 30436 14408 30438
rect 14432 30436 14488 30438
rect 14512 30436 14568 30438
rect 18711 30490 18767 30492
rect 18791 30490 18847 30492
rect 18871 30490 18927 30492
rect 18951 30490 19007 30492
rect 18711 30438 18757 30490
rect 18757 30438 18767 30490
rect 18791 30438 18821 30490
rect 18821 30438 18833 30490
rect 18833 30438 18847 30490
rect 18871 30438 18885 30490
rect 18885 30438 18897 30490
rect 18897 30438 18927 30490
rect 18951 30438 18961 30490
rect 18961 30438 19007 30490
rect 18711 30436 18767 30438
rect 18791 30436 18847 30438
rect 18871 30436 18927 30438
rect 18951 30436 19007 30438
rect 12053 29946 12109 29948
rect 12133 29946 12189 29948
rect 12213 29946 12269 29948
rect 12293 29946 12349 29948
rect 12053 29894 12099 29946
rect 12099 29894 12109 29946
rect 12133 29894 12163 29946
rect 12163 29894 12175 29946
rect 12175 29894 12189 29946
rect 12213 29894 12227 29946
rect 12227 29894 12239 29946
rect 12239 29894 12269 29946
rect 12293 29894 12303 29946
rect 12303 29894 12349 29946
rect 12053 29892 12109 29894
rect 12133 29892 12189 29894
rect 12213 29892 12269 29894
rect 12293 29892 12349 29894
rect 16492 29946 16548 29948
rect 16572 29946 16628 29948
rect 16652 29946 16708 29948
rect 16732 29946 16788 29948
rect 16492 29894 16538 29946
rect 16538 29894 16548 29946
rect 16572 29894 16602 29946
rect 16602 29894 16614 29946
rect 16614 29894 16628 29946
rect 16652 29894 16666 29946
rect 16666 29894 16678 29946
rect 16678 29894 16708 29946
rect 16732 29894 16742 29946
rect 16742 29894 16788 29946
rect 16492 29892 16548 29894
rect 16572 29892 16628 29894
rect 16652 29892 16708 29894
rect 16732 29892 16788 29894
rect 9833 29402 9889 29404
rect 9913 29402 9969 29404
rect 9993 29402 10049 29404
rect 10073 29402 10129 29404
rect 9833 29350 9879 29402
rect 9879 29350 9889 29402
rect 9913 29350 9943 29402
rect 9943 29350 9955 29402
rect 9955 29350 9969 29402
rect 9993 29350 10007 29402
rect 10007 29350 10019 29402
rect 10019 29350 10049 29402
rect 10073 29350 10083 29402
rect 10083 29350 10129 29402
rect 9833 29348 9889 29350
rect 9913 29348 9969 29350
rect 9993 29348 10049 29350
rect 10073 29348 10129 29350
rect 14272 29402 14328 29404
rect 14352 29402 14408 29404
rect 14432 29402 14488 29404
rect 14512 29402 14568 29404
rect 14272 29350 14318 29402
rect 14318 29350 14328 29402
rect 14352 29350 14382 29402
rect 14382 29350 14394 29402
rect 14394 29350 14408 29402
rect 14432 29350 14446 29402
rect 14446 29350 14458 29402
rect 14458 29350 14488 29402
rect 14512 29350 14522 29402
rect 14522 29350 14568 29402
rect 14272 29348 14328 29350
rect 14352 29348 14408 29350
rect 14432 29348 14488 29350
rect 14512 29348 14568 29350
rect 18711 29402 18767 29404
rect 18791 29402 18847 29404
rect 18871 29402 18927 29404
rect 18951 29402 19007 29404
rect 18711 29350 18757 29402
rect 18757 29350 18767 29402
rect 18791 29350 18821 29402
rect 18821 29350 18833 29402
rect 18833 29350 18847 29402
rect 18871 29350 18885 29402
rect 18885 29350 18897 29402
rect 18897 29350 18927 29402
rect 18951 29350 18961 29402
rect 18961 29350 19007 29402
rect 18711 29348 18767 29350
rect 18791 29348 18847 29350
rect 18871 29348 18927 29350
rect 18951 29348 19007 29350
rect 12053 28858 12109 28860
rect 12133 28858 12189 28860
rect 12213 28858 12269 28860
rect 12293 28858 12349 28860
rect 12053 28806 12099 28858
rect 12099 28806 12109 28858
rect 12133 28806 12163 28858
rect 12163 28806 12175 28858
rect 12175 28806 12189 28858
rect 12213 28806 12227 28858
rect 12227 28806 12239 28858
rect 12239 28806 12269 28858
rect 12293 28806 12303 28858
rect 12303 28806 12349 28858
rect 12053 28804 12109 28806
rect 12133 28804 12189 28806
rect 12213 28804 12269 28806
rect 12293 28804 12349 28806
rect 16492 28858 16548 28860
rect 16572 28858 16628 28860
rect 16652 28858 16708 28860
rect 16732 28858 16788 28860
rect 16492 28806 16538 28858
rect 16538 28806 16548 28858
rect 16572 28806 16602 28858
rect 16602 28806 16614 28858
rect 16614 28806 16628 28858
rect 16652 28806 16666 28858
rect 16666 28806 16678 28858
rect 16678 28806 16708 28858
rect 16732 28806 16742 28858
rect 16742 28806 16788 28858
rect 16492 28804 16548 28806
rect 16572 28804 16628 28806
rect 16652 28804 16708 28806
rect 16732 28804 16788 28806
rect 9833 28314 9889 28316
rect 9913 28314 9969 28316
rect 9993 28314 10049 28316
rect 10073 28314 10129 28316
rect 9833 28262 9879 28314
rect 9879 28262 9889 28314
rect 9913 28262 9943 28314
rect 9943 28262 9955 28314
rect 9955 28262 9969 28314
rect 9993 28262 10007 28314
rect 10007 28262 10019 28314
rect 10019 28262 10049 28314
rect 10073 28262 10083 28314
rect 10083 28262 10129 28314
rect 9833 28260 9889 28262
rect 9913 28260 9969 28262
rect 9993 28260 10049 28262
rect 10073 28260 10129 28262
rect 14272 28314 14328 28316
rect 14352 28314 14408 28316
rect 14432 28314 14488 28316
rect 14512 28314 14568 28316
rect 14272 28262 14318 28314
rect 14318 28262 14328 28314
rect 14352 28262 14382 28314
rect 14382 28262 14394 28314
rect 14394 28262 14408 28314
rect 14432 28262 14446 28314
rect 14446 28262 14458 28314
rect 14458 28262 14488 28314
rect 14512 28262 14522 28314
rect 14522 28262 14568 28314
rect 14272 28260 14328 28262
rect 14352 28260 14408 28262
rect 14432 28260 14488 28262
rect 14512 28260 14568 28262
rect 18711 28314 18767 28316
rect 18791 28314 18847 28316
rect 18871 28314 18927 28316
rect 18951 28314 19007 28316
rect 18711 28262 18757 28314
rect 18757 28262 18767 28314
rect 18791 28262 18821 28314
rect 18821 28262 18833 28314
rect 18833 28262 18847 28314
rect 18871 28262 18885 28314
rect 18885 28262 18897 28314
rect 18897 28262 18927 28314
rect 18951 28262 18961 28314
rect 18961 28262 19007 28314
rect 18711 28260 18767 28262
rect 18791 28260 18847 28262
rect 18871 28260 18927 28262
rect 18951 28260 19007 28262
rect 12053 27770 12109 27772
rect 12133 27770 12189 27772
rect 12213 27770 12269 27772
rect 12293 27770 12349 27772
rect 12053 27718 12099 27770
rect 12099 27718 12109 27770
rect 12133 27718 12163 27770
rect 12163 27718 12175 27770
rect 12175 27718 12189 27770
rect 12213 27718 12227 27770
rect 12227 27718 12239 27770
rect 12239 27718 12269 27770
rect 12293 27718 12303 27770
rect 12303 27718 12349 27770
rect 12053 27716 12109 27718
rect 12133 27716 12189 27718
rect 12213 27716 12269 27718
rect 12293 27716 12349 27718
rect 16492 27770 16548 27772
rect 16572 27770 16628 27772
rect 16652 27770 16708 27772
rect 16732 27770 16788 27772
rect 16492 27718 16538 27770
rect 16538 27718 16548 27770
rect 16572 27718 16602 27770
rect 16602 27718 16614 27770
rect 16614 27718 16628 27770
rect 16652 27718 16666 27770
rect 16666 27718 16678 27770
rect 16678 27718 16708 27770
rect 16732 27718 16742 27770
rect 16742 27718 16788 27770
rect 16492 27716 16548 27718
rect 16572 27716 16628 27718
rect 16652 27716 16708 27718
rect 16732 27716 16788 27718
rect 9833 27226 9889 27228
rect 9913 27226 9969 27228
rect 9993 27226 10049 27228
rect 10073 27226 10129 27228
rect 9833 27174 9879 27226
rect 9879 27174 9889 27226
rect 9913 27174 9943 27226
rect 9943 27174 9955 27226
rect 9955 27174 9969 27226
rect 9993 27174 10007 27226
rect 10007 27174 10019 27226
rect 10019 27174 10049 27226
rect 10073 27174 10083 27226
rect 10083 27174 10129 27226
rect 9833 27172 9889 27174
rect 9913 27172 9969 27174
rect 9993 27172 10049 27174
rect 10073 27172 10129 27174
rect 14272 27226 14328 27228
rect 14352 27226 14408 27228
rect 14432 27226 14488 27228
rect 14512 27226 14568 27228
rect 14272 27174 14318 27226
rect 14318 27174 14328 27226
rect 14352 27174 14382 27226
rect 14382 27174 14394 27226
rect 14394 27174 14408 27226
rect 14432 27174 14446 27226
rect 14446 27174 14458 27226
rect 14458 27174 14488 27226
rect 14512 27174 14522 27226
rect 14522 27174 14568 27226
rect 14272 27172 14328 27174
rect 14352 27172 14408 27174
rect 14432 27172 14488 27174
rect 14512 27172 14568 27174
rect 18711 27226 18767 27228
rect 18791 27226 18847 27228
rect 18871 27226 18927 27228
rect 18951 27226 19007 27228
rect 18711 27174 18757 27226
rect 18757 27174 18767 27226
rect 18791 27174 18821 27226
rect 18821 27174 18833 27226
rect 18833 27174 18847 27226
rect 18871 27174 18885 27226
rect 18885 27174 18897 27226
rect 18897 27174 18927 27226
rect 18951 27174 18961 27226
rect 18961 27174 19007 27226
rect 18711 27172 18767 27174
rect 18791 27172 18847 27174
rect 18871 27172 18927 27174
rect 18951 27172 19007 27174
rect 12053 26682 12109 26684
rect 12133 26682 12189 26684
rect 12213 26682 12269 26684
rect 12293 26682 12349 26684
rect 12053 26630 12099 26682
rect 12099 26630 12109 26682
rect 12133 26630 12163 26682
rect 12163 26630 12175 26682
rect 12175 26630 12189 26682
rect 12213 26630 12227 26682
rect 12227 26630 12239 26682
rect 12239 26630 12269 26682
rect 12293 26630 12303 26682
rect 12303 26630 12349 26682
rect 12053 26628 12109 26630
rect 12133 26628 12189 26630
rect 12213 26628 12269 26630
rect 12293 26628 12349 26630
rect 16492 26682 16548 26684
rect 16572 26682 16628 26684
rect 16652 26682 16708 26684
rect 16732 26682 16788 26684
rect 16492 26630 16538 26682
rect 16538 26630 16548 26682
rect 16572 26630 16602 26682
rect 16602 26630 16614 26682
rect 16614 26630 16628 26682
rect 16652 26630 16666 26682
rect 16666 26630 16678 26682
rect 16678 26630 16708 26682
rect 16732 26630 16742 26682
rect 16742 26630 16788 26682
rect 16492 26628 16548 26630
rect 16572 26628 16628 26630
rect 16652 26628 16708 26630
rect 16732 26628 16788 26630
rect 9833 26138 9889 26140
rect 9913 26138 9969 26140
rect 9993 26138 10049 26140
rect 10073 26138 10129 26140
rect 9833 26086 9879 26138
rect 9879 26086 9889 26138
rect 9913 26086 9943 26138
rect 9943 26086 9955 26138
rect 9955 26086 9969 26138
rect 9993 26086 10007 26138
rect 10007 26086 10019 26138
rect 10019 26086 10049 26138
rect 10073 26086 10083 26138
rect 10083 26086 10129 26138
rect 9833 26084 9889 26086
rect 9913 26084 9969 26086
rect 9993 26084 10049 26086
rect 10073 26084 10129 26086
rect 14272 26138 14328 26140
rect 14352 26138 14408 26140
rect 14432 26138 14488 26140
rect 14512 26138 14568 26140
rect 14272 26086 14318 26138
rect 14318 26086 14328 26138
rect 14352 26086 14382 26138
rect 14382 26086 14394 26138
rect 14394 26086 14408 26138
rect 14432 26086 14446 26138
rect 14446 26086 14458 26138
rect 14458 26086 14488 26138
rect 14512 26086 14522 26138
rect 14522 26086 14568 26138
rect 14272 26084 14328 26086
rect 14352 26084 14408 26086
rect 14432 26084 14488 26086
rect 14512 26084 14568 26086
rect 18711 26138 18767 26140
rect 18791 26138 18847 26140
rect 18871 26138 18927 26140
rect 18951 26138 19007 26140
rect 18711 26086 18757 26138
rect 18757 26086 18767 26138
rect 18791 26086 18821 26138
rect 18821 26086 18833 26138
rect 18833 26086 18847 26138
rect 18871 26086 18885 26138
rect 18885 26086 18897 26138
rect 18897 26086 18927 26138
rect 18951 26086 18961 26138
rect 18961 26086 19007 26138
rect 18711 26084 18767 26086
rect 18791 26084 18847 26086
rect 18871 26084 18927 26086
rect 18951 26084 19007 26086
rect 12053 25594 12109 25596
rect 12133 25594 12189 25596
rect 12213 25594 12269 25596
rect 12293 25594 12349 25596
rect 12053 25542 12099 25594
rect 12099 25542 12109 25594
rect 12133 25542 12163 25594
rect 12163 25542 12175 25594
rect 12175 25542 12189 25594
rect 12213 25542 12227 25594
rect 12227 25542 12239 25594
rect 12239 25542 12269 25594
rect 12293 25542 12303 25594
rect 12303 25542 12349 25594
rect 12053 25540 12109 25542
rect 12133 25540 12189 25542
rect 12213 25540 12269 25542
rect 12293 25540 12349 25542
rect 16492 25594 16548 25596
rect 16572 25594 16628 25596
rect 16652 25594 16708 25596
rect 16732 25594 16788 25596
rect 16492 25542 16538 25594
rect 16538 25542 16548 25594
rect 16572 25542 16602 25594
rect 16602 25542 16614 25594
rect 16614 25542 16628 25594
rect 16652 25542 16666 25594
rect 16666 25542 16678 25594
rect 16678 25542 16708 25594
rect 16732 25542 16742 25594
rect 16742 25542 16788 25594
rect 16492 25540 16548 25542
rect 16572 25540 16628 25542
rect 16652 25540 16708 25542
rect 16732 25540 16788 25542
rect 9833 25050 9889 25052
rect 9913 25050 9969 25052
rect 9993 25050 10049 25052
rect 10073 25050 10129 25052
rect 9833 24998 9879 25050
rect 9879 24998 9889 25050
rect 9913 24998 9943 25050
rect 9943 24998 9955 25050
rect 9955 24998 9969 25050
rect 9993 24998 10007 25050
rect 10007 24998 10019 25050
rect 10019 24998 10049 25050
rect 10073 24998 10083 25050
rect 10083 24998 10129 25050
rect 9833 24996 9889 24998
rect 9913 24996 9969 24998
rect 9993 24996 10049 24998
rect 10073 24996 10129 24998
rect 14272 25050 14328 25052
rect 14352 25050 14408 25052
rect 14432 25050 14488 25052
rect 14512 25050 14568 25052
rect 14272 24998 14318 25050
rect 14318 24998 14328 25050
rect 14352 24998 14382 25050
rect 14382 24998 14394 25050
rect 14394 24998 14408 25050
rect 14432 24998 14446 25050
rect 14446 24998 14458 25050
rect 14458 24998 14488 25050
rect 14512 24998 14522 25050
rect 14522 24998 14568 25050
rect 14272 24996 14328 24998
rect 14352 24996 14408 24998
rect 14432 24996 14488 24998
rect 14512 24996 14568 24998
rect 18711 25050 18767 25052
rect 18791 25050 18847 25052
rect 18871 25050 18927 25052
rect 18951 25050 19007 25052
rect 18711 24998 18757 25050
rect 18757 24998 18767 25050
rect 18791 24998 18821 25050
rect 18821 24998 18833 25050
rect 18833 24998 18847 25050
rect 18871 24998 18885 25050
rect 18885 24998 18897 25050
rect 18897 24998 18927 25050
rect 18951 24998 18961 25050
rect 18961 24998 19007 25050
rect 18711 24996 18767 24998
rect 18791 24996 18847 24998
rect 18871 24996 18927 24998
rect 18951 24996 19007 24998
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 12053 24506 12109 24508
rect 12133 24506 12189 24508
rect 12213 24506 12269 24508
rect 12293 24506 12349 24508
rect 12053 24454 12099 24506
rect 12099 24454 12109 24506
rect 12133 24454 12163 24506
rect 12163 24454 12175 24506
rect 12175 24454 12189 24506
rect 12213 24454 12227 24506
rect 12227 24454 12239 24506
rect 12239 24454 12269 24506
rect 12293 24454 12303 24506
rect 12303 24454 12349 24506
rect 12053 24452 12109 24454
rect 12133 24452 12189 24454
rect 12213 24452 12269 24454
rect 12293 24452 12349 24454
rect 16492 24506 16548 24508
rect 16572 24506 16628 24508
rect 16652 24506 16708 24508
rect 16732 24506 16788 24508
rect 16492 24454 16538 24506
rect 16538 24454 16548 24506
rect 16572 24454 16602 24506
rect 16602 24454 16614 24506
rect 16614 24454 16628 24506
rect 16652 24454 16666 24506
rect 16666 24454 16678 24506
rect 16678 24454 16708 24506
rect 16732 24454 16742 24506
rect 16742 24454 16788 24506
rect 16492 24452 16548 24454
rect 16572 24452 16628 24454
rect 16652 24452 16708 24454
rect 16732 24452 16788 24454
rect 9833 23962 9889 23964
rect 9913 23962 9969 23964
rect 9993 23962 10049 23964
rect 10073 23962 10129 23964
rect 9833 23910 9879 23962
rect 9879 23910 9889 23962
rect 9913 23910 9943 23962
rect 9943 23910 9955 23962
rect 9955 23910 9969 23962
rect 9993 23910 10007 23962
rect 10007 23910 10019 23962
rect 10019 23910 10049 23962
rect 10073 23910 10083 23962
rect 10083 23910 10129 23962
rect 9833 23908 9889 23910
rect 9913 23908 9969 23910
rect 9993 23908 10049 23910
rect 10073 23908 10129 23910
rect 14272 23962 14328 23964
rect 14352 23962 14408 23964
rect 14432 23962 14488 23964
rect 14512 23962 14568 23964
rect 14272 23910 14318 23962
rect 14318 23910 14328 23962
rect 14352 23910 14382 23962
rect 14382 23910 14394 23962
rect 14394 23910 14408 23962
rect 14432 23910 14446 23962
rect 14446 23910 14458 23962
rect 14458 23910 14488 23962
rect 14512 23910 14522 23962
rect 14522 23910 14568 23962
rect 14272 23908 14328 23910
rect 14352 23908 14408 23910
rect 14432 23908 14488 23910
rect 14512 23908 14568 23910
rect 18711 23962 18767 23964
rect 18791 23962 18847 23964
rect 18871 23962 18927 23964
rect 18951 23962 19007 23964
rect 18711 23910 18757 23962
rect 18757 23910 18767 23962
rect 18791 23910 18821 23962
rect 18821 23910 18833 23962
rect 18833 23910 18847 23962
rect 18871 23910 18885 23962
rect 18885 23910 18897 23962
rect 18897 23910 18927 23962
rect 18951 23910 18961 23962
rect 18961 23910 19007 23962
rect 18711 23908 18767 23910
rect 18791 23908 18847 23910
rect 18871 23908 18927 23910
rect 18951 23908 19007 23910
rect 12053 23418 12109 23420
rect 12133 23418 12189 23420
rect 12213 23418 12269 23420
rect 12293 23418 12349 23420
rect 12053 23366 12099 23418
rect 12099 23366 12109 23418
rect 12133 23366 12163 23418
rect 12163 23366 12175 23418
rect 12175 23366 12189 23418
rect 12213 23366 12227 23418
rect 12227 23366 12239 23418
rect 12239 23366 12269 23418
rect 12293 23366 12303 23418
rect 12303 23366 12349 23418
rect 12053 23364 12109 23366
rect 12133 23364 12189 23366
rect 12213 23364 12269 23366
rect 12293 23364 12349 23366
rect 16492 23418 16548 23420
rect 16572 23418 16628 23420
rect 16652 23418 16708 23420
rect 16732 23418 16788 23420
rect 16492 23366 16538 23418
rect 16538 23366 16548 23418
rect 16572 23366 16602 23418
rect 16602 23366 16614 23418
rect 16614 23366 16628 23418
rect 16652 23366 16666 23418
rect 16666 23366 16678 23418
rect 16678 23366 16708 23418
rect 16732 23366 16742 23418
rect 16742 23366 16788 23418
rect 16492 23364 16548 23366
rect 16572 23364 16628 23366
rect 16652 23364 16708 23366
rect 16732 23364 16788 23366
rect 9833 22874 9889 22876
rect 9913 22874 9969 22876
rect 9993 22874 10049 22876
rect 10073 22874 10129 22876
rect 9833 22822 9879 22874
rect 9879 22822 9889 22874
rect 9913 22822 9943 22874
rect 9943 22822 9955 22874
rect 9955 22822 9969 22874
rect 9993 22822 10007 22874
rect 10007 22822 10019 22874
rect 10019 22822 10049 22874
rect 10073 22822 10083 22874
rect 10083 22822 10129 22874
rect 9833 22820 9889 22822
rect 9913 22820 9969 22822
rect 9993 22820 10049 22822
rect 10073 22820 10129 22822
rect 14272 22874 14328 22876
rect 14352 22874 14408 22876
rect 14432 22874 14488 22876
rect 14512 22874 14568 22876
rect 14272 22822 14318 22874
rect 14318 22822 14328 22874
rect 14352 22822 14382 22874
rect 14382 22822 14394 22874
rect 14394 22822 14408 22874
rect 14432 22822 14446 22874
rect 14446 22822 14458 22874
rect 14458 22822 14488 22874
rect 14512 22822 14522 22874
rect 14522 22822 14568 22874
rect 14272 22820 14328 22822
rect 14352 22820 14408 22822
rect 14432 22820 14488 22822
rect 14512 22820 14568 22822
rect 18711 22874 18767 22876
rect 18791 22874 18847 22876
rect 18871 22874 18927 22876
rect 18951 22874 19007 22876
rect 18711 22822 18757 22874
rect 18757 22822 18767 22874
rect 18791 22822 18821 22874
rect 18821 22822 18833 22874
rect 18833 22822 18847 22874
rect 18871 22822 18885 22874
rect 18885 22822 18897 22874
rect 18897 22822 18927 22874
rect 18951 22822 18961 22874
rect 18961 22822 19007 22874
rect 18711 22820 18767 22822
rect 18791 22820 18847 22822
rect 18871 22820 18927 22822
rect 18951 22820 19007 22822
rect 12053 22330 12109 22332
rect 12133 22330 12189 22332
rect 12213 22330 12269 22332
rect 12293 22330 12349 22332
rect 12053 22278 12099 22330
rect 12099 22278 12109 22330
rect 12133 22278 12163 22330
rect 12163 22278 12175 22330
rect 12175 22278 12189 22330
rect 12213 22278 12227 22330
rect 12227 22278 12239 22330
rect 12239 22278 12269 22330
rect 12293 22278 12303 22330
rect 12303 22278 12349 22330
rect 12053 22276 12109 22278
rect 12133 22276 12189 22278
rect 12213 22276 12269 22278
rect 12293 22276 12349 22278
rect 16492 22330 16548 22332
rect 16572 22330 16628 22332
rect 16652 22330 16708 22332
rect 16732 22330 16788 22332
rect 16492 22278 16538 22330
rect 16538 22278 16548 22330
rect 16572 22278 16602 22330
rect 16602 22278 16614 22330
rect 16614 22278 16628 22330
rect 16652 22278 16666 22330
rect 16666 22278 16678 22330
rect 16678 22278 16708 22330
rect 16732 22278 16742 22330
rect 16742 22278 16788 22330
rect 16492 22276 16548 22278
rect 16572 22276 16628 22278
rect 16652 22276 16708 22278
rect 16732 22276 16788 22278
rect 9833 21786 9889 21788
rect 9913 21786 9969 21788
rect 9993 21786 10049 21788
rect 10073 21786 10129 21788
rect 9833 21734 9879 21786
rect 9879 21734 9889 21786
rect 9913 21734 9943 21786
rect 9943 21734 9955 21786
rect 9955 21734 9969 21786
rect 9993 21734 10007 21786
rect 10007 21734 10019 21786
rect 10019 21734 10049 21786
rect 10073 21734 10083 21786
rect 10083 21734 10129 21786
rect 9833 21732 9889 21734
rect 9913 21732 9969 21734
rect 9993 21732 10049 21734
rect 10073 21732 10129 21734
rect 14272 21786 14328 21788
rect 14352 21786 14408 21788
rect 14432 21786 14488 21788
rect 14512 21786 14568 21788
rect 14272 21734 14318 21786
rect 14318 21734 14328 21786
rect 14352 21734 14382 21786
rect 14382 21734 14394 21786
rect 14394 21734 14408 21786
rect 14432 21734 14446 21786
rect 14446 21734 14458 21786
rect 14458 21734 14488 21786
rect 14512 21734 14522 21786
rect 14522 21734 14568 21786
rect 14272 21732 14328 21734
rect 14352 21732 14408 21734
rect 14432 21732 14488 21734
rect 14512 21732 14568 21734
rect 18711 21786 18767 21788
rect 18791 21786 18847 21788
rect 18871 21786 18927 21788
rect 18951 21786 19007 21788
rect 18711 21734 18757 21786
rect 18757 21734 18767 21786
rect 18791 21734 18821 21786
rect 18821 21734 18833 21786
rect 18833 21734 18847 21786
rect 18871 21734 18885 21786
rect 18885 21734 18897 21786
rect 18897 21734 18927 21786
rect 18951 21734 18961 21786
rect 18961 21734 19007 21786
rect 18711 21732 18767 21734
rect 18791 21732 18847 21734
rect 18871 21732 18927 21734
rect 18951 21732 19007 21734
rect 12053 21242 12109 21244
rect 12133 21242 12189 21244
rect 12213 21242 12269 21244
rect 12293 21242 12349 21244
rect 12053 21190 12099 21242
rect 12099 21190 12109 21242
rect 12133 21190 12163 21242
rect 12163 21190 12175 21242
rect 12175 21190 12189 21242
rect 12213 21190 12227 21242
rect 12227 21190 12239 21242
rect 12239 21190 12269 21242
rect 12293 21190 12303 21242
rect 12303 21190 12349 21242
rect 12053 21188 12109 21190
rect 12133 21188 12189 21190
rect 12213 21188 12269 21190
rect 12293 21188 12349 21190
rect 16492 21242 16548 21244
rect 16572 21242 16628 21244
rect 16652 21242 16708 21244
rect 16732 21242 16788 21244
rect 16492 21190 16538 21242
rect 16538 21190 16548 21242
rect 16572 21190 16602 21242
rect 16602 21190 16614 21242
rect 16614 21190 16628 21242
rect 16652 21190 16666 21242
rect 16666 21190 16678 21242
rect 16678 21190 16708 21242
rect 16732 21190 16742 21242
rect 16742 21190 16788 21242
rect 16492 21188 16548 21190
rect 16572 21188 16628 21190
rect 16652 21188 16708 21190
rect 16732 21188 16788 21190
rect 9833 20698 9889 20700
rect 9913 20698 9969 20700
rect 9993 20698 10049 20700
rect 10073 20698 10129 20700
rect 9833 20646 9879 20698
rect 9879 20646 9889 20698
rect 9913 20646 9943 20698
rect 9943 20646 9955 20698
rect 9955 20646 9969 20698
rect 9993 20646 10007 20698
rect 10007 20646 10019 20698
rect 10019 20646 10049 20698
rect 10073 20646 10083 20698
rect 10083 20646 10129 20698
rect 9833 20644 9889 20646
rect 9913 20644 9969 20646
rect 9993 20644 10049 20646
rect 10073 20644 10129 20646
rect 14272 20698 14328 20700
rect 14352 20698 14408 20700
rect 14432 20698 14488 20700
rect 14512 20698 14568 20700
rect 14272 20646 14318 20698
rect 14318 20646 14328 20698
rect 14352 20646 14382 20698
rect 14382 20646 14394 20698
rect 14394 20646 14408 20698
rect 14432 20646 14446 20698
rect 14446 20646 14458 20698
rect 14458 20646 14488 20698
rect 14512 20646 14522 20698
rect 14522 20646 14568 20698
rect 14272 20644 14328 20646
rect 14352 20644 14408 20646
rect 14432 20644 14488 20646
rect 14512 20644 14568 20646
rect 18711 20698 18767 20700
rect 18791 20698 18847 20700
rect 18871 20698 18927 20700
rect 18951 20698 19007 20700
rect 18711 20646 18757 20698
rect 18757 20646 18767 20698
rect 18791 20646 18821 20698
rect 18821 20646 18833 20698
rect 18833 20646 18847 20698
rect 18871 20646 18885 20698
rect 18885 20646 18897 20698
rect 18897 20646 18927 20698
rect 18951 20646 18961 20698
rect 18961 20646 19007 20698
rect 18711 20644 18767 20646
rect 18791 20644 18847 20646
rect 18871 20644 18927 20646
rect 18951 20644 19007 20646
rect 12053 20154 12109 20156
rect 12133 20154 12189 20156
rect 12213 20154 12269 20156
rect 12293 20154 12349 20156
rect 12053 20102 12099 20154
rect 12099 20102 12109 20154
rect 12133 20102 12163 20154
rect 12163 20102 12175 20154
rect 12175 20102 12189 20154
rect 12213 20102 12227 20154
rect 12227 20102 12239 20154
rect 12239 20102 12269 20154
rect 12293 20102 12303 20154
rect 12303 20102 12349 20154
rect 12053 20100 12109 20102
rect 12133 20100 12189 20102
rect 12213 20100 12269 20102
rect 12293 20100 12349 20102
rect 16492 20154 16548 20156
rect 16572 20154 16628 20156
rect 16652 20154 16708 20156
rect 16732 20154 16788 20156
rect 16492 20102 16538 20154
rect 16538 20102 16548 20154
rect 16572 20102 16602 20154
rect 16602 20102 16614 20154
rect 16614 20102 16628 20154
rect 16652 20102 16666 20154
rect 16666 20102 16678 20154
rect 16678 20102 16708 20154
rect 16732 20102 16742 20154
rect 16742 20102 16788 20154
rect 16492 20100 16548 20102
rect 16572 20100 16628 20102
rect 16652 20100 16708 20102
rect 16732 20100 16788 20102
rect 9833 19610 9889 19612
rect 9913 19610 9969 19612
rect 9993 19610 10049 19612
rect 10073 19610 10129 19612
rect 9833 19558 9879 19610
rect 9879 19558 9889 19610
rect 9913 19558 9943 19610
rect 9943 19558 9955 19610
rect 9955 19558 9969 19610
rect 9993 19558 10007 19610
rect 10007 19558 10019 19610
rect 10019 19558 10049 19610
rect 10073 19558 10083 19610
rect 10083 19558 10129 19610
rect 9833 19556 9889 19558
rect 9913 19556 9969 19558
rect 9993 19556 10049 19558
rect 10073 19556 10129 19558
rect 14272 19610 14328 19612
rect 14352 19610 14408 19612
rect 14432 19610 14488 19612
rect 14512 19610 14568 19612
rect 14272 19558 14318 19610
rect 14318 19558 14328 19610
rect 14352 19558 14382 19610
rect 14382 19558 14394 19610
rect 14394 19558 14408 19610
rect 14432 19558 14446 19610
rect 14446 19558 14458 19610
rect 14458 19558 14488 19610
rect 14512 19558 14522 19610
rect 14522 19558 14568 19610
rect 14272 19556 14328 19558
rect 14352 19556 14408 19558
rect 14432 19556 14488 19558
rect 14512 19556 14568 19558
rect 18711 19610 18767 19612
rect 18791 19610 18847 19612
rect 18871 19610 18927 19612
rect 18951 19610 19007 19612
rect 18711 19558 18757 19610
rect 18757 19558 18767 19610
rect 18791 19558 18821 19610
rect 18821 19558 18833 19610
rect 18833 19558 18847 19610
rect 18871 19558 18885 19610
rect 18885 19558 18897 19610
rect 18897 19558 18927 19610
rect 18951 19558 18961 19610
rect 18961 19558 19007 19610
rect 18711 19556 18767 19558
rect 18791 19556 18847 19558
rect 18871 19556 18927 19558
rect 18951 19556 19007 19558
rect 12053 19066 12109 19068
rect 12133 19066 12189 19068
rect 12213 19066 12269 19068
rect 12293 19066 12349 19068
rect 12053 19014 12099 19066
rect 12099 19014 12109 19066
rect 12133 19014 12163 19066
rect 12163 19014 12175 19066
rect 12175 19014 12189 19066
rect 12213 19014 12227 19066
rect 12227 19014 12239 19066
rect 12239 19014 12269 19066
rect 12293 19014 12303 19066
rect 12303 19014 12349 19066
rect 12053 19012 12109 19014
rect 12133 19012 12189 19014
rect 12213 19012 12269 19014
rect 12293 19012 12349 19014
rect 16492 19066 16548 19068
rect 16572 19066 16628 19068
rect 16652 19066 16708 19068
rect 16732 19066 16788 19068
rect 16492 19014 16538 19066
rect 16538 19014 16548 19066
rect 16572 19014 16602 19066
rect 16602 19014 16614 19066
rect 16614 19014 16628 19066
rect 16652 19014 16666 19066
rect 16666 19014 16678 19066
rect 16678 19014 16708 19066
rect 16732 19014 16742 19066
rect 16742 19014 16788 19066
rect 16492 19012 16548 19014
rect 16572 19012 16628 19014
rect 16652 19012 16708 19014
rect 16732 19012 16788 19014
rect 9833 18522 9889 18524
rect 9913 18522 9969 18524
rect 9993 18522 10049 18524
rect 10073 18522 10129 18524
rect 9833 18470 9879 18522
rect 9879 18470 9889 18522
rect 9913 18470 9943 18522
rect 9943 18470 9955 18522
rect 9955 18470 9969 18522
rect 9993 18470 10007 18522
rect 10007 18470 10019 18522
rect 10019 18470 10049 18522
rect 10073 18470 10083 18522
rect 10083 18470 10129 18522
rect 9833 18468 9889 18470
rect 9913 18468 9969 18470
rect 9993 18468 10049 18470
rect 10073 18468 10129 18470
rect 14272 18522 14328 18524
rect 14352 18522 14408 18524
rect 14432 18522 14488 18524
rect 14512 18522 14568 18524
rect 14272 18470 14318 18522
rect 14318 18470 14328 18522
rect 14352 18470 14382 18522
rect 14382 18470 14394 18522
rect 14394 18470 14408 18522
rect 14432 18470 14446 18522
rect 14446 18470 14458 18522
rect 14458 18470 14488 18522
rect 14512 18470 14522 18522
rect 14522 18470 14568 18522
rect 14272 18468 14328 18470
rect 14352 18468 14408 18470
rect 14432 18468 14488 18470
rect 14512 18468 14568 18470
rect 18711 18522 18767 18524
rect 18791 18522 18847 18524
rect 18871 18522 18927 18524
rect 18951 18522 19007 18524
rect 18711 18470 18757 18522
rect 18757 18470 18767 18522
rect 18791 18470 18821 18522
rect 18821 18470 18833 18522
rect 18833 18470 18847 18522
rect 18871 18470 18885 18522
rect 18885 18470 18897 18522
rect 18897 18470 18927 18522
rect 18951 18470 18961 18522
rect 18961 18470 19007 18522
rect 18711 18468 18767 18470
rect 18791 18468 18847 18470
rect 18871 18468 18927 18470
rect 18951 18468 19007 18470
rect 12053 17978 12109 17980
rect 12133 17978 12189 17980
rect 12213 17978 12269 17980
rect 12293 17978 12349 17980
rect 12053 17926 12099 17978
rect 12099 17926 12109 17978
rect 12133 17926 12163 17978
rect 12163 17926 12175 17978
rect 12175 17926 12189 17978
rect 12213 17926 12227 17978
rect 12227 17926 12239 17978
rect 12239 17926 12269 17978
rect 12293 17926 12303 17978
rect 12303 17926 12349 17978
rect 12053 17924 12109 17926
rect 12133 17924 12189 17926
rect 12213 17924 12269 17926
rect 12293 17924 12349 17926
rect 16492 17978 16548 17980
rect 16572 17978 16628 17980
rect 16652 17978 16708 17980
rect 16732 17978 16788 17980
rect 16492 17926 16538 17978
rect 16538 17926 16548 17978
rect 16572 17926 16602 17978
rect 16602 17926 16614 17978
rect 16614 17926 16628 17978
rect 16652 17926 16666 17978
rect 16666 17926 16678 17978
rect 16678 17926 16708 17978
rect 16732 17926 16742 17978
rect 16742 17926 16788 17978
rect 16492 17924 16548 17926
rect 16572 17924 16628 17926
rect 16652 17924 16708 17926
rect 16732 17924 16788 17926
rect 9833 17434 9889 17436
rect 9913 17434 9969 17436
rect 9993 17434 10049 17436
rect 10073 17434 10129 17436
rect 9833 17382 9879 17434
rect 9879 17382 9889 17434
rect 9913 17382 9943 17434
rect 9943 17382 9955 17434
rect 9955 17382 9969 17434
rect 9993 17382 10007 17434
rect 10007 17382 10019 17434
rect 10019 17382 10049 17434
rect 10073 17382 10083 17434
rect 10083 17382 10129 17434
rect 9833 17380 9889 17382
rect 9913 17380 9969 17382
rect 9993 17380 10049 17382
rect 10073 17380 10129 17382
rect 14272 17434 14328 17436
rect 14352 17434 14408 17436
rect 14432 17434 14488 17436
rect 14512 17434 14568 17436
rect 14272 17382 14318 17434
rect 14318 17382 14328 17434
rect 14352 17382 14382 17434
rect 14382 17382 14394 17434
rect 14394 17382 14408 17434
rect 14432 17382 14446 17434
rect 14446 17382 14458 17434
rect 14458 17382 14488 17434
rect 14512 17382 14522 17434
rect 14522 17382 14568 17434
rect 14272 17380 14328 17382
rect 14352 17380 14408 17382
rect 14432 17380 14488 17382
rect 14512 17380 14568 17382
rect 18711 17434 18767 17436
rect 18791 17434 18847 17436
rect 18871 17434 18927 17436
rect 18951 17434 19007 17436
rect 18711 17382 18757 17434
rect 18757 17382 18767 17434
rect 18791 17382 18821 17434
rect 18821 17382 18833 17434
rect 18833 17382 18847 17434
rect 18871 17382 18885 17434
rect 18885 17382 18897 17434
rect 18897 17382 18927 17434
rect 18951 17382 18961 17434
rect 18961 17382 19007 17434
rect 18711 17380 18767 17382
rect 18791 17380 18847 17382
rect 18871 17380 18927 17382
rect 18951 17380 19007 17382
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 9833 16346 9889 16348
rect 9913 16346 9969 16348
rect 9993 16346 10049 16348
rect 10073 16346 10129 16348
rect 9833 16294 9879 16346
rect 9879 16294 9889 16346
rect 9913 16294 9943 16346
rect 9943 16294 9955 16346
rect 9955 16294 9969 16346
rect 9993 16294 10007 16346
rect 10007 16294 10019 16346
rect 10019 16294 10049 16346
rect 10073 16294 10083 16346
rect 10083 16294 10129 16346
rect 9833 16292 9889 16294
rect 9913 16292 9969 16294
rect 9993 16292 10049 16294
rect 10073 16292 10129 16294
rect 14272 16346 14328 16348
rect 14352 16346 14408 16348
rect 14432 16346 14488 16348
rect 14512 16346 14568 16348
rect 14272 16294 14318 16346
rect 14318 16294 14328 16346
rect 14352 16294 14382 16346
rect 14382 16294 14394 16346
rect 14394 16294 14408 16346
rect 14432 16294 14446 16346
rect 14446 16294 14458 16346
rect 14458 16294 14488 16346
rect 14512 16294 14522 16346
rect 14522 16294 14568 16346
rect 14272 16292 14328 16294
rect 14352 16292 14408 16294
rect 14432 16292 14488 16294
rect 14512 16292 14568 16294
rect 18711 16346 18767 16348
rect 18791 16346 18847 16348
rect 18871 16346 18927 16348
rect 18951 16346 19007 16348
rect 18711 16294 18757 16346
rect 18757 16294 18767 16346
rect 18791 16294 18821 16346
rect 18821 16294 18833 16346
rect 18833 16294 18847 16346
rect 18871 16294 18885 16346
rect 18885 16294 18897 16346
rect 18897 16294 18927 16346
rect 18951 16294 18961 16346
rect 18961 16294 19007 16346
rect 18711 16292 18767 16294
rect 18791 16292 18847 16294
rect 18871 16292 18927 16294
rect 18951 16292 19007 16294
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 9833 15258 9889 15260
rect 9913 15258 9969 15260
rect 9993 15258 10049 15260
rect 10073 15258 10129 15260
rect 9833 15206 9879 15258
rect 9879 15206 9889 15258
rect 9913 15206 9943 15258
rect 9943 15206 9955 15258
rect 9955 15206 9969 15258
rect 9993 15206 10007 15258
rect 10007 15206 10019 15258
rect 10019 15206 10049 15258
rect 10073 15206 10083 15258
rect 10083 15206 10129 15258
rect 9833 15204 9889 15206
rect 9913 15204 9969 15206
rect 9993 15204 10049 15206
rect 10073 15204 10129 15206
rect 14272 15258 14328 15260
rect 14352 15258 14408 15260
rect 14432 15258 14488 15260
rect 14512 15258 14568 15260
rect 14272 15206 14318 15258
rect 14318 15206 14328 15258
rect 14352 15206 14382 15258
rect 14382 15206 14394 15258
rect 14394 15206 14408 15258
rect 14432 15206 14446 15258
rect 14446 15206 14458 15258
rect 14458 15206 14488 15258
rect 14512 15206 14522 15258
rect 14522 15206 14568 15258
rect 14272 15204 14328 15206
rect 14352 15204 14408 15206
rect 14432 15204 14488 15206
rect 14512 15204 14568 15206
rect 18711 15258 18767 15260
rect 18791 15258 18847 15260
rect 18871 15258 18927 15260
rect 18951 15258 19007 15260
rect 18711 15206 18757 15258
rect 18757 15206 18767 15258
rect 18791 15206 18821 15258
rect 18821 15206 18833 15258
rect 18833 15206 18847 15258
rect 18871 15206 18885 15258
rect 18885 15206 18897 15258
rect 18897 15206 18927 15258
rect 18951 15206 18961 15258
rect 18961 15206 19007 15258
rect 18711 15204 18767 15206
rect 18791 15204 18847 15206
rect 18871 15204 18927 15206
rect 18951 15204 19007 15206
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 9833 14170 9889 14172
rect 9913 14170 9969 14172
rect 9993 14170 10049 14172
rect 10073 14170 10129 14172
rect 9833 14118 9879 14170
rect 9879 14118 9889 14170
rect 9913 14118 9943 14170
rect 9943 14118 9955 14170
rect 9955 14118 9969 14170
rect 9993 14118 10007 14170
rect 10007 14118 10019 14170
rect 10019 14118 10049 14170
rect 10073 14118 10083 14170
rect 10083 14118 10129 14170
rect 9833 14116 9889 14118
rect 9913 14116 9969 14118
rect 9993 14116 10049 14118
rect 10073 14116 10129 14118
rect 14272 14170 14328 14172
rect 14352 14170 14408 14172
rect 14432 14170 14488 14172
rect 14512 14170 14568 14172
rect 14272 14118 14318 14170
rect 14318 14118 14328 14170
rect 14352 14118 14382 14170
rect 14382 14118 14394 14170
rect 14394 14118 14408 14170
rect 14432 14118 14446 14170
rect 14446 14118 14458 14170
rect 14458 14118 14488 14170
rect 14512 14118 14522 14170
rect 14522 14118 14568 14170
rect 14272 14116 14328 14118
rect 14352 14116 14408 14118
rect 14432 14116 14488 14118
rect 14512 14116 14568 14118
rect 18711 14170 18767 14172
rect 18791 14170 18847 14172
rect 18871 14170 18927 14172
rect 18951 14170 19007 14172
rect 18711 14118 18757 14170
rect 18757 14118 18767 14170
rect 18791 14118 18821 14170
rect 18821 14118 18833 14170
rect 18833 14118 18847 14170
rect 18871 14118 18885 14170
rect 18885 14118 18897 14170
rect 18897 14118 18927 14170
rect 18951 14118 18961 14170
rect 18961 14118 19007 14170
rect 18711 14116 18767 14118
rect 18791 14116 18847 14118
rect 18871 14116 18927 14118
rect 18951 14116 19007 14118
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 9833 13082 9889 13084
rect 9913 13082 9969 13084
rect 9993 13082 10049 13084
rect 10073 13082 10129 13084
rect 9833 13030 9879 13082
rect 9879 13030 9889 13082
rect 9913 13030 9943 13082
rect 9943 13030 9955 13082
rect 9955 13030 9969 13082
rect 9993 13030 10007 13082
rect 10007 13030 10019 13082
rect 10019 13030 10049 13082
rect 10073 13030 10083 13082
rect 10083 13030 10129 13082
rect 9833 13028 9889 13030
rect 9913 13028 9969 13030
rect 9993 13028 10049 13030
rect 10073 13028 10129 13030
rect 14272 13082 14328 13084
rect 14352 13082 14408 13084
rect 14432 13082 14488 13084
rect 14512 13082 14568 13084
rect 14272 13030 14318 13082
rect 14318 13030 14328 13082
rect 14352 13030 14382 13082
rect 14382 13030 14394 13082
rect 14394 13030 14408 13082
rect 14432 13030 14446 13082
rect 14446 13030 14458 13082
rect 14458 13030 14488 13082
rect 14512 13030 14522 13082
rect 14522 13030 14568 13082
rect 14272 13028 14328 13030
rect 14352 13028 14408 13030
rect 14432 13028 14488 13030
rect 14512 13028 14568 13030
rect 18711 13082 18767 13084
rect 18791 13082 18847 13084
rect 18871 13082 18927 13084
rect 18951 13082 19007 13084
rect 18711 13030 18757 13082
rect 18757 13030 18767 13082
rect 18791 13030 18821 13082
rect 18821 13030 18833 13082
rect 18833 13030 18847 13082
rect 18871 13030 18885 13082
rect 18885 13030 18897 13082
rect 18897 13030 18927 13082
rect 18951 13030 18961 13082
rect 18961 13030 19007 13082
rect 18711 13028 18767 13030
rect 18791 13028 18847 13030
rect 18871 13028 18927 13030
rect 18951 13028 19007 13030
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 9833 11994 9889 11996
rect 9913 11994 9969 11996
rect 9993 11994 10049 11996
rect 10073 11994 10129 11996
rect 9833 11942 9879 11994
rect 9879 11942 9889 11994
rect 9913 11942 9943 11994
rect 9943 11942 9955 11994
rect 9955 11942 9969 11994
rect 9993 11942 10007 11994
rect 10007 11942 10019 11994
rect 10019 11942 10049 11994
rect 10073 11942 10083 11994
rect 10083 11942 10129 11994
rect 9833 11940 9889 11942
rect 9913 11940 9969 11942
rect 9993 11940 10049 11942
rect 10073 11940 10129 11942
rect 14272 11994 14328 11996
rect 14352 11994 14408 11996
rect 14432 11994 14488 11996
rect 14512 11994 14568 11996
rect 14272 11942 14318 11994
rect 14318 11942 14328 11994
rect 14352 11942 14382 11994
rect 14382 11942 14394 11994
rect 14394 11942 14408 11994
rect 14432 11942 14446 11994
rect 14446 11942 14458 11994
rect 14458 11942 14488 11994
rect 14512 11942 14522 11994
rect 14522 11942 14568 11994
rect 14272 11940 14328 11942
rect 14352 11940 14408 11942
rect 14432 11940 14488 11942
rect 14512 11940 14568 11942
rect 18711 11994 18767 11996
rect 18791 11994 18847 11996
rect 18871 11994 18927 11996
rect 18951 11994 19007 11996
rect 18711 11942 18757 11994
rect 18757 11942 18767 11994
rect 18791 11942 18821 11994
rect 18821 11942 18833 11994
rect 18833 11942 18847 11994
rect 18871 11942 18885 11994
rect 18885 11942 18897 11994
rect 18897 11942 18927 11994
rect 18951 11942 18961 11994
rect 18961 11942 19007 11994
rect 18711 11940 18767 11942
rect 18791 11940 18847 11942
rect 18871 11940 18927 11942
rect 18951 11940 19007 11942
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 9833 10906 9889 10908
rect 9913 10906 9969 10908
rect 9993 10906 10049 10908
rect 10073 10906 10129 10908
rect 9833 10854 9879 10906
rect 9879 10854 9889 10906
rect 9913 10854 9943 10906
rect 9943 10854 9955 10906
rect 9955 10854 9969 10906
rect 9993 10854 10007 10906
rect 10007 10854 10019 10906
rect 10019 10854 10049 10906
rect 10073 10854 10083 10906
rect 10083 10854 10129 10906
rect 9833 10852 9889 10854
rect 9913 10852 9969 10854
rect 9993 10852 10049 10854
rect 10073 10852 10129 10854
rect 14272 10906 14328 10908
rect 14352 10906 14408 10908
rect 14432 10906 14488 10908
rect 14512 10906 14568 10908
rect 14272 10854 14318 10906
rect 14318 10854 14328 10906
rect 14352 10854 14382 10906
rect 14382 10854 14394 10906
rect 14394 10854 14408 10906
rect 14432 10854 14446 10906
rect 14446 10854 14458 10906
rect 14458 10854 14488 10906
rect 14512 10854 14522 10906
rect 14522 10854 14568 10906
rect 14272 10852 14328 10854
rect 14352 10852 14408 10854
rect 14432 10852 14488 10854
rect 14512 10852 14568 10854
rect 18711 10906 18767 10908
rect 18791 10906 18847 10908
rect 18871 10906 18927 10908
rect 18951 10906 19007 10908
rect 18711 10854 18757 10906
rect 18757 10854 18767 10906
rect 18791 10854 18821 10906
rect 18821 10854 18833 10906
rect 18833 10854 18847 10906
rect 18871 10854 18885 10906
rect 18885 10854 18897 10906
rect 18897 10854 18927 10906
rect 18951 10854 18961 10906
rect 18961 10854 19007 10906
rect 18711 10852 18767 10854
rect 18791 10852 18847 10854
rect 18871 10852 18927 10854
rect 18951 10852 19007 10854
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 9833 9818 9889 9820
rect 9913 9818 9969 9820
rect 9993 9818 10049 9820
rect 10073 9818 10129 9820
rect 9833 9766 9879 9818
rect 9879 9766 9889 9818
rect 9913 9766 9943 9818
rect 9943 9766 9955 9818
rect 9955 9766 9969 9818
rect 9993 9766 10007 9818
rect 10007 9766 10019 9818
rect 10019 9766 10049 9818
rect 10073 9766 10083 9818
rect 10083 9766 10129 9818
rect 9833 9764 9889 9766
rect 9913 9764 9969 9766
rect 9993 9764 10049 9766
rect 10073 9764 10129 9766
rect 14272 9818 14328 9820
rect 14352 9818 14408 9820
rect 14432 9818 14488 9820
rect 14512 9818 14568 9820
rect 14272 9766 14318 9818
rect 14318 9766 14328 9818
rect 14352 9766 14382 9818
rect 14382 9766 14394 9818
rect 14394 9766 14408 9818
rect 14432 9766 14446 9818
rect 14446 9766 14458 9818
rect 14458 9766 14488 9818
rect 14512 9766 14522 9818
rect 14522 9766 14568 9818
rect 14272 9764 14328 9766
rect 14352 9764 14408 9766
rect 14432 9764 14488 9766
rect 14512 9764 14568 9766
rect 18711 9818 18767 9820
rect 18791 9818 18847 9820
rect 18871 9818 18927 9820
rect 18951 9818 19007 9820
rect 18711 9766 18757 9818
rect 18757 9766 18767 9818
rect 18791 9766 18821 9818
rect 18821 9766 18833 9818
rect 18833 9766 18847 9818
rect 18871 9766 18885 9818
rect 18885 9766 18897 9818
rect 18897 9766 18927 9818
rect 18951 9766 18961 9818
rect 18961 9766 19007 9818
rect 18711 9764 18767 9766
rect 18791 9764 18847 9766
rect 18871 9764 18927 9766
rect 18951 9764 19007 9766
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 9833 8730 9889 8732
rect 9913 8730 9969 8732
rect 9993 8730 10049 8732
rect 10073 8730 10129 8732
rect 9833 8678 9879 8730
rect 9879 8678 9889 8730
rect 9913 8678 9943 8730
rect 9943 8678 9955 8730
rect 9955 8678 9969 8730
rect 9993 8678 10007 8730
rect 10007 8678 10019 8730
rect 10019 8678 10049 8730
rect 10073 8678 10083 8730
rect 10083 8678 10129 8730
rect 9833 8676 9889 8678
rect 9913 8676 9969 8678
rect 9993 8676 10049 8678
rect 10073 8676 10129 8678
rect 14272 8730 14328 8732
rect 14352 8730 14408 8732
rect 14432 8730 14488 8732
rect 14512 8730 14568 8732
rect 14272 8678 14318 8730
rect 14318 8678 14328 8730
rect 14352 8678 14382 8730
rect 14382 8678 14394 8730
rect 14394 8678 14408 8730
rect 14432 8678 14446 8730
rect 14446 8678 14458 8730
rect 14458 8678 14488 8730
rect 14512 8678 14522 8730
rect 14522 8678 14568 8730
rect 14272 8676 14328 8678
rect 14352 8676 14408 8678
rect 14432 8676 14488 8678
rect 14512 8676 14568 8678
rect 18711 8730 18767 8732
rect 18791 8730 18847 8732
rect 18871 8730 18927 8732
rect 18951 8730 19007 8732
rect 18711 8678 18757 8730
rect 18757 8678 18767 8730
rect 18791 8678 18821 8730
rect 18821 8678 18833 8730
rect 18833 8678 18847 8730
rect 18871 8678 18885 8730
rect 18885 8678 18897 8730
rect 18897 8678 18927 8730
rect 18951 8678 18961 8730
rect 18961 8678 19007 8730
rect 18711 8676 18767 8678
rect 18791 8676 18847 8678
rect 18871 8676 18927 8678
rect 18951 8676 19007 8678
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
<< metal3 >>
rect 0 47970 800 48000
rect 933 47970 999 47973
rect 0 47968 999 47970
rect 0 47912 938 47968
rect 994 47912 999 47968
rect 0 47910 999 47912
rect 0 47880 800 47910
rect 933 47907 999 47910
rect 3165 47360 3481 47361
rect 3165 47296 3171 47360
rect 3235 47296 3251 47360
rect 3315 47296 3331 47360
rect 3395 47296 3411 47360
rect 3475 47296 3481 47360
rect 3165 47295 3481 47296
rect 7604 47360 7920 47361
rect 7604 47296 7610 47360
rect 7674 47296 7690 47360
rect 7754 47296 7770 47360
rect 7834 47296 7850 47360
rect 7914 47296 7920 47360
rect 7604 47295 7920 47296
rect 12043 47360 12359 47361
rect 12043 47296 12049 47360
rect 12113 47296 12129 47360
rect 12193 47296 12209 47360
rect 12273 47296 12289 47360
rect 12353 47296 12359 47360
rect 12043 47295 12359 47296
rect 16482 47360 16798 47361
rect 16482 47296 16488 47360
rect 16552 47296 16568 47360
rect 16632 47296 16648 47360
rect 16712 47296 16728 47360
rect 16792 47296 16798 47360
rect 16482 47295 16798 47296
rect 5384 46816 5700 46817
rect 5384 46752 5390 46816
rect 5454 46752 5470 46816
rect 5534 46752 5550 46816
rect 5614 46752 5630 46816
rect 5694 46752 5700 46816
rect 5384 46751 5700 46752
rect 9823 46816 10139 46817
rect 9823 46752 9829 46816
rect 9893 46752 9909 46816
rect 9973 46752 9989 46816
rect 10053 46752 10069 46816
rect 10133 46752 10139 46816
rect 9823 46751 10139 46752
rect 14262 46816 14578 46817
rect 14262 46752 14268 46816
rect 14332 46752 14348 46816
rect 14412 46752 14428 46816
rect 14492 46752 14508 46816
rect 14572 46752 14578 46816
rect 14262 46751 14578 46752
rect 18701 46816 19017 46817
rect 18701 46752 18707 46816
rect 18771 46752 18787 46816
rect 18851 46752 18867 46816
rect 18931 46752 18947 46816
rect 19011 46752 19017 46816
rect 18701 46751 19017 46752
rect 3165 46272 3481 46273
rect 3165 46208 3171 46272
rect 3235 46208 3251 46272
rect 3315 46208 3331 46272
rect 3395 46208 3411 46272
rect 3475 46208 3481 46272
rect 3165 46207 3481 46208
rect 7604 46272 7920 46273
rect 7604 46208 7610 46272
rect 7674 46208 7690 46272
rect 7754 46208 7770 46272
rect 7834 46208 7850 46272
rect 7914 46208 7920 46272
rect 7604 46207 7920 46208
rect 12043 46272 12359 46273
rect 12043 46208 12049 46272
rect 12113 46208 12129 46272
rect 12193 46208 12209 46272
rect 12273 46208 12289 46272
rect 12353 46208 12359 46272
rect 12043 46207 12359 46208
rect 16482 46272 16798 46273
rect 16482 46208 16488 46272
rect 16552 46208 16568 46272
rect 16632 46208 16648 46272
rect 16712 46208 16728 46272
rect 16792 46208 16798 46272
rect 16482 46207 16798 46208
rect 5384 45728 5700 45729
rect 5384 45664 5390 45728
rect 5454 45664 5470 45728
rect 5534 45664 5550 45728
rect 5614 45664 5630 45728
rect 5694 45664 5700 45728
rect 5384 45663 5700 45664
rect 9823 45728 10139 45729
rect 9823 45664 9829 45728
rect 9893 45664 9909 45728
rect 9973 45664 9989 45728
rect 10053 45664 10069 45728
rect 10133 45664 10139 45728
rect 9823 45663 10139 45664
rect 14262 45728 14578 45729
rect 14262 45664 14268 45728
rect 14332 45664 14348 45728
rect 14412 45664 14428 45728
rect 14492 45664 14508 45728
rect 14572 45664 14578 45728
rect 14262 45663 14578 45664
rect 18701 45728 19017 45729
rect 18701 45664 18707 45728
rect 18771 45664 18787 45728
rect 18851 45664 18867 45728
rect 18931 45664 18947 45728
rect 19011 45664 19017 45728
rect 18701 45663 19017 45664
rect 3165 45184 3481 45185
rect 3165 45120 3171 45184
rect 3235 45120 3251 45184
rect 3315 45120 3331 45184
rect 3395 45120 3411 45184
rect 3475 45120 3481 45184
rect 3165 45119 3481 45120
rect 7604 45184 7920 45185
rect 7604 45120 7610 45184
rect 7674 45120 7690 45184
rect 7754 45120 7770 45184
rect 7834 45120 7850 45184
rect 7914 45120 7920 45184
rect 7604 45119 7920 45120
rect 12043 45184 12359 45185
rect 12043 45120 12049 45184
rect 12113 45120 12129 45184
rect 12193 45120 12209 45184
rect 12273 45120 12289 45184
rect 12353 45120 12359 45184
rect 12043 45119 12359 45120
rect 16482 45184 16798 45185
rect 16482 45120 16488 45184
rect 16552 45120 16568 45184
rect 16632 45120 16648 45184
rect 16712 45120 16728 45184
rect 16792 45120 16798 45184
rect 16482 45119 16798 45120
rect 5384 44640 5700 44641
rect 5384 44576 5390 44640
rect 5454 44576 5470 44640
rect 5534 44576 5550 44640
rect 5614 44576 5630 44640
rect 5694 44576 5700 44640
rect 5384 44575 5700 44576
rect 9823 44640 10139 44641
rect 9823 44576 9829 44640
rect 9893 44576 9909 44640
rect 9973 44576 9989 44640
rect 10053 44576 10069 44640
rect 10133 44576 10139 44640
rect 9823 44575 10139 44576
rect 14262 44640 14578 44641
rect 14262 44576 14268 44640
rect 14332 44576 14348 44640
rect 14412 44576 14428 44640
rect 14492 44576 14508 44640
rect 14572 44576 14578 44640
rect 14262 44575 14578 44576
rect 18701 44640 19017 44641
rect 18701 44576 18707 44640
rect 18771 44576 18787 44640
rect 18851 44576 18867 44640
rect 18931 44576 18947 44640
rect 19011 44576 19017 44640
rect 18701 44575 19017 44576
rect 0 44434 800 44464
rect 933 44434 999 44437
rect 0 44432 999 44434
rect 0 44376 938 44432
rect 994 44376 999 44432
rect 0 44374 999 44376
rect 0 44344 800 44374
rect 933 44371 999 44374
rect 3165 44096 3481 44097
rect 3165 44032 3171 44096
rect 3235 44032 3251 44096
rect 3315 44032 3331 44096
rect 3395 44032 3411 44096
rect 3475 44032 3481 44096
rect 3165 44031 3481 44032
rect 7604 44096 7920 44097
rect 7604 44032 7610 44096
rect 7674 44032 7690 44096
rect 7754 44032 7770 44096
rect 7834 44032 7850 44096
rect 7914 44032 7920 44096
rect 7604 44031 7920 44032
rect 12043 44096 12359 44097
rect 12043 44032 12049 44096
rect 12113 44032 12129 44096
rect 12193 44032 12209 44096
rect 12273 44032 12289 44096
rect 12353 44032 12359 44096
rect 12043 44031 12359 44032
rect 16482 44096 16798 44097
rect 16482 44032 16488 44096
rect 16552 44032 16568 44096
rect 16632 44032 16648 44096
rect 16712 44032 16728 44096
rect 16792 44032 16798 44096
rect 16482 44031 16798 44032
rect 5384 43552 5700 43553
rect 5384 43488 5390 43552
rect 5454 43488 5470 43552
rect 5534 43488 5550 43552
rect 5614 43488 5630 43552
rect 5694 43488 5700 43552
rect 5384 43487 5700 43488
rect 9823 43552 10139 43553
rect 9823 43488 9829 43552
rect 9893 43488 9909 43552
rect 9973 43488 9989 43552
rect 10053 43488 10069 43552
rect 10133 43488 10139 43552
rect 9823 43487 10139 43488
rect 14262 43552 14578 43553
rect 14262 43488 14268 43552
rect 14332 43488 14348 43552
rect 14412 43488 14428 43552
rect 14492 43488 14508 43552
rect 14572 43488 14578 43552
rect 14262 43487 14578 43488
rect 18701 43552 19017 43553
rect 18701 43488 18707 43552
rect 18771 43488 18787 43552
rect 18851 43488 18867 43552
rect 18931 43488 18947 43552
rect 19011 43488 19017 43552
rect 18701 43487 19017 43488
rect 3165 43008 3481 43009
rect 3165 42944 3171 43008
rect 3235 42944 3251 43008
rect 3315 42944 3331 43008
rect 3395 42944 3411 43008
rect 3475 42944 3481 43008
rect 3165 42943 3481 42944
rect 7604 43008 7920 43009
rect 7604 42944 7610 43008
rect 7674 42944 7690 43008
rect 7754 42944 7770 43008
rect 7834 42944 7850 43008
rect 7914 42944 7920 43008
rect 7604 42943 7920 42944
rect 12043 43008 12359 43009
rect 12043 42944 12049 43008
rect 12113 42944 12129 43008
rect 12193 42944 12209 43008
rect 12273 42944 12289 43008
rect 12353 42944 12359 43008
rect 12043 42943 12359 42944
rect 16482 43008 16798 43009
rect 16482 42944 16488 43008
rect 16552 42944 16568 43008
rect 16632 42944 16648 43008
rect 16712 42944 16728 43008
rect 16792 42944 16798 43008
rect 16482 42943 16798 42944
rect 5384 42464 5700 42465
rect 5384 42400 5390 42464
rect 5454 42400 5470 42464
rect 5534 42400 5550 42464
rect 5614 42400 5630 42464
rect 5694 42400 5700 42464
rect 5384 42399 5700 42400
rect 9823 42464 10139 42465
rect 9823 42400 9829 42464
rect 9893 42400 9909 42464
rect 9973 42400 9989 42464
rect 10053 42400 10069 42464
rect 10133 42400 10139 42464
rect 9823 42399 10139 42400
rect 14262 42464 14578 42465
rect 14262 42400 14268 42464
rect 14332 42400 14348 42464
rect 14412 42400 14428 42464
rect 14492 42400 14508 42464
rect 14572 42400 14578 42464
rect 14262 42399 14578 42400
rect 18701 42464 19017 42465
rect 18701 42400 18707 42464
rect 18771 42400 18787 42464
rect 18851 42400 18867 42464
rect 18931 42400 18947 42464
rect 19011 42400 19017 42464
rect 18701 42399 19017 42400
rect 3165 41920 3481 41921
rect 3165 41856 3171 41920
rect 3235 41856 3251 41920
rect 3315 41856 3331 41920
rect 3395 41856 3411 41920
rect 3475 41856 3481 41920
rect 3165 41855 3481 41856
rect 7604 41920 7920 41921
rect 7604 41856 7610 41920
rect 7674 41856 7690 41920
rect 7754 41856 7770 41920
rect 7834 41856 7850 41920
rect 7914 41856 7920 41920
rect 7604 41855 7920 41856
rect 12043 41920 12359 41921
rect 12043 41856 12049 41920
rect 12113 41856 12129 41920
rect 12193 41856 12209 41920
rect 12273 41856 12289 41920
rect 12353 41856 12359 41920
rect 12043 41855 12359 41856
rect 16482 41920 16798 41921
rect 16482 41856 16488 41920
rect 16552 41856 16568 41920
rect 16632 41856 16648 41920
rect 16712 41856 16728 41920
rect 16792 41856 16798 41920
rect 16482 41855 16798 41856
rect 5384 41376 5700 41377
rect 5384 41312 5390 41376
rect 5454 41312 5470 41376
rect 5534 41312 5550 41376
rect 5614 41312 5630 41376
rect 5694 41312 5700 41376
rect 5384 41311 5700 41312
rect 9823 41376 10139 41377
rect 9823 41312 9829 41376
rect 9893 41312 9909 41376
rect 9973 41312 9989 41376
rect 10053 41312 10069 41376
rect 10133 41312 10139 41376
rect 9823 41311 10139 41312
rect 14262 41376 14578 41377
rect 14262 41312 14268 41376
rect 14332 41312 14348 41376
rect 14412 41312 14428 41376
rect 14492 41312 14508 41376
rect 14572 41312 14578 41376
rect 14262 41311 14578 41312
rect 18701 41376 19017 41377
rect 18701 41312 18707 41376
rect 18771 41312 18787 41376
rect 18851 41312 18867 41376
rect 18931 41312 18947 41376
rect 19011 41312 19017 41376
rect 18701 41311 19017 41312
rect 0 40898 800 40928
rect 933 40898 999 40901
rect 0 40896 999 40898
rect 0 40840 938 40896
rect 994 40840 999 40896
rect 0 40838 999 40840
rect 0 40808 800 40838
rect 933 40835 999 40838
rect 3165 40832 3481 40833
rect 3165 40768 3171 40832
rect 3235 40768 3251 40832
rect 3315 40768 3331 40832
rect 3395 40768 3411 40832
rect 3475 40768 3481 40832
rect 3165 40767 3481 40768
rect 7604 40832 7920 40833
rect 7604 40768 7610 40832
rect 7674 40768 7690 40832
rect 7754 40768 7770 40832
rect 7834 40768 7850 40832
rect 7914 40768 7920 40832
rect 7604 40767 7920 40768
rect 12043 40832 12359 40833
rect 12043 40768 12049 40832
rect 12113 40768 12129 40832
rect 12193 40768 12209 40832
rect 12273 40768 12289 40832
rect 12353 40768 12359 40832
rect 12043 40767 12359 40768
rect 16482 40832 16798 40833
rect 16482 40768 16488 40832
rect 16552 40768 16568 40832
rect 16632 40768 16648 40832
rect 16712 40768 16728 40832
rect 16792 40768 16798 40832
rect 16482 40767 16798 40768
rect 5384 40288 5700 40289
rect 5384 40224 5390 40288
rect 5454 40224 5470 40288
rect 5534 40224 5550 40288
rect 5614 40224 5630 40288
rect 5694 40224 5700 40288
rect 5384 40223 5700 40224
rect 9823 40288 10139 40289
rect 9823 40224 9829 40288
rect 9893 40224 9909 40288
rect 9973 40224 9989 40288
rect 10053 40224 10069 40288
rect 10133 40224 10139 40288
rect 9823 40223 10139 40224
rect 14262 40288 14578 40289
rect 14262 40224 14268 40288
rect 14332 40224 14348 40288
rect 14412 40224 14428 40288
rect 14492 40224 14508 40288
rect 14572 40224 14578 40288
rect 14262 40223 14578 40224
rect 18701 40288 19017 40289
rect 18701 40224 18707 40288
rect 18771 40224 18787 40288
rect 18851 40224 18867 40288
rect 18931 40224 18947 40288
rect 19011 40224 19017 40288
rect 18701 40223 19017 40224
rect 3165 39744 3481 39745
rect 3165 39680 3171 39744
rect 3235 39680 3251 39744
rect 3315 39680 3331 39744
rect 3395 39680 3411 39744
rect 3475 39680 3481 39744
rect 3165 39679 3481 39680
rect 7604 39744 7920 39745
rect 7604 39680 7610 39744
rect 7674 39680 7690 39744
rect 7754 39680 7770 39744
rect 7834 39680 7850 39744
rect 7914 39680 7920 39744
rect 7604 39679 7920 39680
rect 12043 39744 12359 39745
rect 12043 39680 12049 39744
rect 12113 39680 12129 39744
rect 12193 39680 12209 39744
rect 12273 39680 12289 39744
rect 12353 39680 12359 39744
rect 12043 39679 12359 39680
rect 16482 39744 16798 39745
rect 16482 39680 16488 39744
rect 16552 39680 16568 39744
rect 16632 39680 16648 39744
rect 16712 39680 16728 39744
rect 16792 39680 16798 39744
rect 16482 39679 16798 39680
rect 5384 39200 5700 39201
rect 5384 39136 5390 39200
rect 5454 39136 5470 39200
rect 5534 39136 5550 39200
rect 5614 39136 5630 39200
rect 5694 39136 5700 39200
rect 5384 39135 5700 39136
rect 9823 39200 10139 39201
rect 9823 39136 9829 39200
rect 9893 39136 9909 39200
rect 9973 39136 9989 39200
rect 10053 39136 10069 39200
rect 10133 39136 10139 39200
rect 9823 39135 10139 39136
rect 14262 39200 14578 39201
rect 14262 39136 14268 39200
rect 14332 39136 14348 39200
rect 14412 39136 14428 39200
rect 14492 39136 14508 39200
rect 14572 39136 14578 39200
rect 14262 39135 14578 39136
rect 18701 39200 19017 39201
rect 18701 39136 18707 39200
rect 18771 39136 18787 39200
rect 18851 39136 18867 39200
rect 18931 39136 18947 39200
rect 19011 39136 19017 39200
rect 18701 39135 19017 39136
rect 3165 38656 3481 38657
rect 3165 38592 3171 38656
rect 3235 38592 3251 38656
rect 3315 38592 3331 38656
rect 3395 38592 3411 38656
rect 3475 38592 3481 38656
rect 3165 38591 3481 38592
rect 7604 38656 7920 38657
rect 7604 38592 7610 38656
rect 7674 38592 7690 38656
rect 7754 38592 7770 38656
rect 7834 38592 7850 38656
rect 7914 38592 7920 38656
rect 7604 38591 7920 38592
rect 12043 38656 12359 38657
rect 12043 38592 12049 38656
rect 12113 38592 12129 38656
rect 12193 38592 12209 38656
rect 12273 38592 12289 38656
rect 12353 38592 12359 38656
rect 12043 38591 12359 38592
rect 16482 38656 16798 38657
rect 16482 38592 16488 38656
rect 16552 38592 16568 38656
rect 16632 38592 16648 38656
rect 16712 38592 16728 38656
rect 16792 38592 16798 38656
rect 16482 38591 16798 38592
rect 5384 38112 5700 38113
rect 5384 38048 5390 38112
rect 5454 38048 5470 38112
rect 5534 38048 5550 38112
rect 5614 38048 5630 38112
rect 5694 38048 5700 38112
rect 5384 38047 5700 38048
rect 9823 38112 10139 38113
rect 9823 38048 9829 38112
rect 9893 38048 9909 38112
rect 9973 38048 9989 38112
rect 10053 38048 10069 38112
rect 10133 38048 10139 38112
rect 9823 38047 10139 38048
rect 14262 38112 14578 38113
rect 14262 38048 14268 38112
rect 14332 38048 14348 38112
rect 14412 38048 14428 38112
rect 14492 38048 14508 38112
rect 14572 38048 14578 38112
rect 14262 38047 14578 38048
rect 18701 38112 19017 38113
rect 18701 38048 18707 38112
rect 18771 38048 18787 38112
rect 18851 38048 18867 38112
rect 18931 38048 18947 38112
rect 19011 38048 19017 38112
rect 18701 38047 19017 38048
rect 3165 37568 3481 37569
rect 3165 37504 3171 37568
rect 3235 37504 3251 37568
rect 3315 37504 3331 37568
rect 3395 37504 3411 37568
rect 3475 37504 3481 37568
rect 3165 37503 3481 37504
rect 7604 37568 7920 37569
rect 7604 37504 7610 37568
rect 7674 37504 7690 37568
rect 7754 37504 7770 37568
rect 7834 37504 7850 37568
rect 7914 37504 7920 37568
rect 7604 37503 7920 37504
rect 12043 37568 12359 37569
rect 12043 37504 12049 37568
rect 12113 37504 12129 37568
rect 12193 37504 12209 37568
rect 12273 37504 12289 37568
rect 12353 37504 12359 37568
rect 12043 37503 12359 37504
rect 16482 37568 16798 37569
rect 16482 37504 16488 37568
rect 16552 37504 16568 37568
rect 16632 37504 16648 37568
rect 16712 37504 16728 37568
rect 16792 37504 16798 37568
rect 16482 37503 16798 37504
rect 0 37362 800 37392
rect 933 37362 999 37365
rect 0 37360 999 37362
rect 0 37304 938 37360
rect 994 37304 999 37360
rect 0 37302 999 37304
rect 0 37272 800 37302
rect 933 37299 999 37302
rect 5384 37024 5700 37025
rect 5384 36960 5390 37024
rect 5454 36960 5470 37024
rect 5534 36960 5550 37024
rect 5614 36960 5630 37024
rect 5694 36960 5700 37024
rect 5384 36959 5700 36960
rect 9823 37024 10139 37025
rect 9823 36960 9829 37024
rect 9893 36960 9909 37024
rect 9973 36960 9989 37024
rect 10053 36960 10069 37024
rect 10133 36960 10139 37024
rect 9823 36959 10139 36960
rect 14262 37024 14578 37025
rect 14262 36960 14268 37024
rect 14332 36960 14348 37024
rect 14412 36960 14428 37024
rect 14492 36960 14508 37024
rect 14572 36960 14578 37024
rect 14262 36959 14578 36960
rect 18701 37024 19017 37025
rect 18701 36960 18707 37024
rect 18771 36960 18787 37024
rect 18851 36960 18867 37024
rect 18931 36960 18947 37024
rect 19011 36960 19017 37024
rect 18701 36959 19017 36960
rect 3165 36480 3481 36481
rect 3165 36416 3171 36480
rect 3235 36416 3251 36480
rect 3315 36416 3331 36480
rect 3395 36416 3411 36480
rect 3475 36416 3481 36480
rect 3165 36415 3481 36416
rect 7604 36480 7920 36481
rect 7604 36416 7610 36480
rect 7674 36416 7690 36480
rect 7754 36416 7770 36480
rect 7834 36416 7850 36480
rect 7914 36416 7920 36480
rect 7604 36415 7920 36416
rect 12043 36480 12359 36481
rect 12043 36416 12049 36480
rect 12113 36416 12129 36480
rect 12193 36416 12209 36480
rect 12273 36416 12289 36480
rect 12353 36416 12359 36480
rect 12043 36415 12359 36416
rect 16482 36480 16798 36481
rect 16482 36416 16488 36480
rect 16552 36416 16568 36480
rect 16632 36416 16648 36480
rect 16712 36416 16728 36480
rect 16792 36416 16798 36480
rect 16482 36415 16798 36416
rect 5384 35936 5700 35937
rect 5384 35872 5390 35936
rect 5454 35872 5470 35936
rect 5534 35872 5550 35936
rect 5614 35872 5630 35936
rect 5694 35872 5700 35936
rect 5384 35871 5700 35872
rect 9823 35936 10139 35937
rect 9823 35872 9829 35936
rect 9893 35872 9909 35936
rect 9973 35872 9989 35936
rect 10053 35872 10069 35936
rect 10133 35872 10139 35936
rect 9823 35871 10139 35872
rect 14262 35936 14578 35937
rect 14262 35872 14268 35936
rect 14332 35872 14348 35936
rect 14412 35872 14428 35936
rect 14492 35872 14508 35936
rect 14572 35872 14578 35936
rect 14262 35871 14578 35872
rect 18701 35936 19017 35937
rect 18701 35872 18707 35936
rect 18771 35872 18787 35936
rect 18851 35872 18867 35936
rect 18931 35872 18947 35936
rect 19011 35872 19017 35936
rect 18701 35871 19017 35872
rect 3165 35392 3481 35393
rect 3165 35328 3171 35392
rect 3235 35328 3251 35392
rect 3315 35328 3331 35392
rect 3395 35328 3411 35392
rect 3475 35328 3481 35392
rect 3165 35327 3481 35328
rect 7604 35392 7920 35393
rect 7604 35328 7610 35392
rect 7674 35328 7690 35392
rect 7754 35328 7770 35392
rect 7834 35328 7850 35392
rect 7914 35328 7920 35392
rect 7604 35327 7920 35328
rect 12043 35392 12359 35393
rect 12043 35328 12049 35392
rect 12113 35328 12129 35392
rect 12193 35328 12209 35392
rect 12273 35328 12289 35392
rect 12353 35328 12359 35392
rect 12043 35327 12359 35328
rect 16482 35392 16798 35393
rect 16482 35328 16488 35392
rect 16552 35328 16568 35392
rect 16632 35328 16648 35392
rect 16712 35328 16728 35392
rect 16792 35328 16798 35392
rect 16482 35327 16798 35328
rect 5384 34848 5700 34849
rect 5384 34784 5390 34848
rect 5454 34784 5470 34848
rect 5534 34784 5550 34848
rect 5614 34784 5630 34848
rect 5694 34784 5700 34848
rect 5384 34783 5700 34784
rect 9823 34848 10139 34849
rect 9823 34784 9829 34848
rect 9893 34784 9909 34848
rect 9973 34784 9989 34848
rect 10053 34784 10069 34848
rect 10133 34784 10139 34848
rect 9823 34783 10139 34784
rect 14262 34848 14578 34849
rect 14262 34784 14268 34848
rect 14332 34784 14348 34848
rect 14412 34784 14428 34848
rect 14492 34784 14508 34848
rect 14572 34784 14578 34848
rect 14262 34783 14578 34784
rect 18701 34848 19017 34849
rect 18701 34784 18707 34848
rect 18771 34784 18787 34848
rect 18851 34784 18867 34848
rect 18931 34784 18947 34848
rect 19011 34784 19017 34848
rect 18701 34783 19017 34784
rect 3165 34304 3481 34305
rect 3165 34240 3171 34304
rect 3235 34240 3251 34304
rect 3315 34240 3331 34304
rect 3395 34240 3411 34304
rect 3475 34240 3481 34304
rect 3165 34239 3481 34240
rect 7604 34304 7920 34305
rect 7604 34240 7610 34304
rect 7674 34240 7690 34304
rect 7754 34240 7770 34304
rect 7834 34240 7850 34304
rect 7914 34240 7920 34304
rect 7604 34239 7920 34240
rect 12043 34304 12359 34305
rect 12043 34240 12049 34304
rect 12113 34240 12129 34304
rect 12193 34240 12209 34304
rect 12273 34240 12289 34304
rect 12353 34240 12359 34304
rect 12043 34239 12359 34240
rect 16482 34304 16798 34305
rect 16482 34240 16488 34304
rect 16552 34240 16568 34304
rect 16632 34240 16648 34304
rect 16712 34240 16728 34304
rect 16792 34240 16798 34304
rect 16482 34239 16798 34240
rect 0 33826 800 33856
rect 933 33826 999 33829
rect 0 33824 999 33826
rect 0 33768 938 33824
rect 994 33768 999 33824
rect 0 33766 999 33768
rect 0 33736 800 33766
rect 933 33763 999 33766
rect 5384 33760 5700 33761
rect 5384 33696 5390 33760
rect 5454 33696 5470 33760
rect 5534 33696 5550 33760
rect 5614 33696 5630 33760
rect 5694 33696 5700 33760
rect 5384 33695 5700 33696
rect 9823 33760 10139 33761
rect 9823 33696 9829 33760
rect 9893 33696 9909 33760
rect 9973 33696 9989 33760
rect 10053 33696 10069 33760
rect 10133 33696 10139 33760
rect 9823 33695 10139 33696
rect 14262 33760 14578 33761
rect 14262 33696 14268 33760
rect 14332 33696 14348 33760
rect 14412 33696 14428 33760
rect 14492 33696 14508 33760
rect 14572 33696 14578 33760
rect 14262 33695 14578 33696
rect 18701 33760 19017 33761
rect 18701 33696 18707 33760
rect 18771 33696 18787 33760
rect 18851 33696 18867 33760
rect 18931 33696 18947 33760
rect 19011 33696 19017 33760
rect 18701 33695 19017 33696
rect 3165 33216 3481 33217
rect 3165 33152 3171 33216
rect 3235 33152 3251 33216
rect 3315 33152 3331 33216
rect 3395 33152 3411 33216
rect 3475 33152 3481 33216
rect 3165 33151 3481 33152
rect 7604 33216 7920 33217
rect 7604 33152 7610 33216
rect 7674 33152 7690 33216
rect 7754 33152 7770 33216
rect 7834 33152 7850 33216
rect 7914 33152 7920 33216
rect 7604 33151 7920 33152
rect 12043 33216 12359 33217
rect 12043 33152 12049 33216
rect 12113 33152 12129 33216
rect 12193 33152 12209 33216
rect 12273 33152 12289 33216
rect 12353 33152 12359 33216
rect 12043 33151 12359 33152
rect 16482 33216 16798 33217
rect 16482 33152 16488 33216
rect 16552 33152 16568 33216
rect 16632 33152 16648 33216
rect 16712 33152 16728 33216
rect 16792 33152 16798 33216
rect 16482 33151 16798 33152
rect 5384 32672 5700 32673
rect 5384 32608 5390 32672
rect 5454 32608 5470 32672
rect 5534 32608 5550 32672
rect 5614 32608 5630 32672
rect 5694 32608 5700 32672
rect 5384 32607 5700 32608
rect 9823 32672 10139 32673
rect 9823 32608 9829 32672
rect 9893 32608 9909 32672
rect 9973 32608 9989 32672
rect 10053 32608 10069 32672
rect 10133 32608 10139 32672
rect 9823 32607 10139 32608
rect 14262 32672 14578 32673
rect 14262 32608 14268 32672
rect 14332 32608 14348 32672
rect 14412 32608 14428 32672
rect 14492 32608 14508 32672
rect 14572 32608 14578 32672
rect 14262 32607 14578 32608
rect 18701 32672 19017 32673
rect 18701 32608 18707 32672
rect 18771 32608 18787 32672
rect 18851 32608 18867 32672
rect 18931 32608 18947 32672
rect 19011 32608 19017 32672
rect 18701 32607 19017 32608
rect 3165 32128 3481 32129
rect 3165 32064 3171 32128
rect 3235 32064 3251 32128
rect 3315 32064 3331 32128
rect 3395 32064 3411 32128
rect 3475 32064 3481 32128
rect 3165 32063 3481 32064
rect 7604 32128 7920 32129
rect 7604 32064 7610 32128
rect 7674 32064 7690 32128
rect 7754 32064 7770 32128
rect 7834 32064 7850 32128
rect 7914 32064 7920 32128
rect 7604 32063 7920 32064
rect 12043 32128 12359 32129
rect 12043 32064 12049 32128
rect 12113 32064 12129 32128
rect 12193 32064 12209 32128
rect 12273 32064 12289 32128
rect 12353 32064 12359 32128
rect 12043 32063 12359 32064
rect 16482 32128 16798 32129
rect 16482 32064 16488 32128
rect 16552 32064 16568 32128
rect 16632 32064 16648 32128
rect 16712 32064 16728 32128
rect 16792 32064 16798 32128
rect 16482 32063 16798 32064
rect 5384 31584 5700 31585
rect 5384 31520 5390 31584
rect 5454 31520 5470 31584
rect 5534 31520 5550 31584
rect 5614 31520 5630 31584
rect 5694 31520 5700 31584
rect 5384 31519 5700 31520
rect 9823 31584 10139 31585
rect 9823 31520 9829 31584
rect 9893 31520 9909 31584
rect 9973 31520 9989 31584
rect 10053 31520 10069 31584
rect 10133 31520 10139 31584
rect 9823 31519 10139 31520
rect 14262 31584 14578 31585
rect 14262 31520 14268 31584
rect 14332 31520 14348 31584
rect 14412 31520 14428 31584
rect 14492 31520 14508 31584
rect 14572 31520 14578 31584
rect 14262 31519 14578 31520
rect 18701 31584 19017 31585
rect 18701 31520 18707 31584
rect 18771 31520 18787 31584
rect 18851 31520 18867 31584
rect 18931 31520 18947 31584
rect 19011 31520 19017 31584
rect 18701 31519 19017 31520
rect 3165 31040 3481 31041
rect 3165 30976 3171 31040
rect 3235 30976 3251 31040
rect 3315 30976 3331 31040
rect 3395 30976 3411 31040
rect 3475 30976 3481 31040
rect 3165 30975 3481 30976
rect 7604 31040 7920 31041
rect 7604 30976 7610 31040
rect 7674 30976 7690 31040
rect 7754 30976 7770 31040
rect 7834 30976 7850 31040
rect 7914 30976 7920 31040
rect 7604 30975 7920 30976
rect 12043 31040 12359 31041
rect 12043 30976 12049 31040
rect 12113 30976 12129 31040
rect 12193 30976 12209 31040
rect 12273 30976 12289 31040
rect 12353 30976 12359 31040
rect 12043 30975 12359 30976
rect 16482 31040 16798 31041
rect 16482 30976 16488 31040
rect 16552 30976 16568 31040
rect 16632 30976 16648 31040
rect 16712 30976 16728 31040
rect 16792 30976 16798 31040
rect 16482 30975 16798 30976
rect 5384 30496 5700 30497
rect 5384 30432 5390 30496
rect 5454 30432 5470 30496
rect 5534 30432 5550 30496
rect 5614 30432 5630 30496
rect 5694 30432 5700 30496
rect 5384 30431 5700 30432
rect 9823 30496 10139 30497
rect 9823 30432 9829 30496
rect 9893 30432 9909 30496
rect 9973 30432 9989 30496
rect 10053 30432 10069 30496
rect 10133 30432 10139 30496
rect 9823 30431 10139 30432
rect 14262 30496 14578 30497
rect 14262 30432 14268 30496
rect 14332 30432 14348 30496
rect 14412 30432 14428 30496
rect 14492 30432 14508 30496
rect 14572 30432 14578 30496
rect 14262 30431 14578 30432
rect 18701 30496 19017 30497
rect 18701 30432 18707 30496
rect 18771 30432 18787 30496
rect 18851 30432 18867 30496
rect 18931 30432 18947 30496
rect 19011 30432 19017 30496
rect 18701 30431 19017 30432
rect 4705 30428 4771 30429
rect 4654 30426 4660 30428
rect 4614 30366 4660 30426
rect 4724 30424 4771 30428
rect 4766 30368 4771 30424
rect 4654 30364 4660 30366
rect 4724 30364 4771 30368
rect 4705 30363 4771 30364
rect 0 30290 800 30320
rect 933 30290 999 30293
rect 0 30288 999 30290
rect 0 30232 938 30288
rect 994 30232 999 30288
rect 0 30230 999 30232
rect 0 30200 800 30230
rect 933 30227 999 30230
rect 3165 29952 3481 29953
rect 3165 29888 3171 29952
rect 3235 29888 3251 29952
rect 3315 29888 3331 29952
rect 3395 29888 3411 29952
rect 3475 29888 3481 29952
rect 3165 29887 3481 29888
rect 7604 29952 7920 29953
rect 7604 29888 7610 29952
rect 7674 29888 7690 29952
rect 7754 29888 7770 29952
rect 7834 29888 7850 29952
rect 7914 29888 7920 29952
rect 7604 29887 7920 29888
rect 12043 29952 12359 29953
rect 12043 29888 12049 29952
rect 12113 29888 12129 29952
rect 12193 29888 12209 29952
rect 12273 29888 12289 29952
rect 12353 29888 12359 29952
rect 12043 29887 12359 29888
rect 16482 29952 16798 29953
rect 16482 29888 16488 29952
rect 16552 29888 16568 29952
rect 16632 29888 16648 29952
rect 16712 29888 16728 29952
rect 16792 29888 16798 29952
rect 16482 29887 16798 29888
rect 5384 29408 5700 29409
rect 5384 29344 5390 29408
rect 5454 29344 5470 29408
rect 5534 29344 5550 29408
rect 5614 29344 5630 29408
rect 5694 29344 5700 29408
rect 5384 29343 5700 29344
rect 9823 29408 10139 29409
rect 9823 29344 9829 29408
rect 9893 29344 9909 29408
rect 9973 29344 9989 29408
rect 10053 29344 10069 29408
rect 10133 29344 10139 29408
rect 9823 29343 10139 29344
rect 14262 29408 14578 29409
rect 14262 29344 14268 29408
rect 14332 29344 14348 29408
rect 14412 29344 14428 29408
rect 14492 29344 14508 29408
rect 14572 29344 14578 29408
rect 14262 29343 14578 29344
rect 18701 29408 19017 29409
rect 18701 29344 18707 29408
rect 18771 29344 18787 29408
rect 18851 29344 18867 29408
rect 18931 29344 18947 29408
rect 19011 29344 19017 29408
rect 18701 29343 19017 29344
rect 8109 29068 8175 29069
rect 8109 29064 8156 29068
rect 8220 29066 8226 29068
rect 8109 29008 8114 29064
rect 8109 29004 8156 29008
rect 8220 29006 8266 29066
rect 8220 29004 8226 29006
rect 8109 29003 8175 29004
rect 3165 28864 3481 28865
rect 3165 28800 3171 28864
rect 3235 28800 3251 28864
rect 3315 28800 3331 28864
rect 3395 28800 3411 28864
rect 3475 28800 3481 28864
rect 3165 28799 3481 28800
rect 7604 28864 7920 28865
rect 7604 28800 7610 28864
rect 7674 28800 7690 28864
rect 7754 28800 7770 28864
rect 7834 28800 7850 28864
rect 7914 28800 7920 28864
rect 7604 28799 7920 28800
rect 12043 28864 12359 28865
rect 12043 28800 12049 28864
rect 12113 28800 12129 28864
rect 12193 28800 12209 28864
rect 12273 28800 12289 28864
rect 12353 28800 12359 28864
rect 12043 28799 12359 28800
rect 16482 28864 16798 28865
rect 16482 28800 16488 28864
rect 16552 28800 16568 28864
rect 16632 28800 16648 28864
rect 16712 28800 16728 28864
rect 16792 28800 16798 28864
rect 16482 28799 16798 28800
rect 5384 28320 5700 28321
rect 5384 28256 5390 28320
rect 5454 28256 5470 28320
rect 5534 28256 5550 28320
rect 5614 28256 5630 28320
rect 5694 28256 5700 28320
rect 5384 28255 5700 28256
rect 9823 28320 10139 28321
rect 9823 28256 9829 28320
rect 9893 28256 9909 28320
rect 9973 28256 9989 28320
rect 10053 28256 10069 28320
rect 10133 28256 10139 28320
rect 9823 28255 10139 28256
rect 14262 28320 14578 28321
rect 14262 28256 14268 28320
rect 14332 28256 14348 28320
rect 14412 28256 14428 28320
rect 14492 28256 14508 28320
rect 14572 28256 14578 28320
rect 14262 28255 14578 28256
rect 18701 28320 19017 28321
rect 18701 28256 18707 28320
rect 18771 28256 18787 28320
rect 18851 28256 18867 28320
rect 18931 28256 18947 28320
rect 19011 28256 19017 28320
rect 18701 28255 19017 28256
rect 3165 27776 3481 27777
rect 3165 27712 3171 27776
rect 3235 27712 3251 27776
rect 3315 27712 3331 27776
rect 3395 27712 3411 27776
rect 3475 27712 3481 27776
rect 3165 27711 3481 27712
rect 7604 27776 7920 27777
rect 7604 27712 7610 27776
rect 7674 27712 7690 27776
rect 7754 27712 7770 27776
rect 7834 27712 7850 27776
rect 7914 27712 7920 27776
rect 7604 27711 7920 27712
rect 12043 27776 12359 27777
rect 12043 27712 12049 27776
rect 12113 27712 12129 27776
rect 12193 27712 12209 27776
rect 12273 27712 12289 27776
rect 12353 27712 12359 27776
rect 12043 27711 12359 27712
rect 16482 27776 16798 27777
rect 16482 27712 16488 27776
rect 16552 27712 16568 27776
rect 16632 27712 16648 27776
rect 16712 27712 16728 27776
rect 16792 27712 16798 27776
rect 16482 27711 16798 27712
rect 4245 27708 4311 27709
rect 4245 27704 4292 27708
rect 4356 27706 4362 27708
rect 4245 27648 4250 27704
rect 4245 27644 4292 27648
rect 4356 27646 4402 27706
rect 4356 27644 4362 27646
rect 4245 27643 4311 27644
rect 5384 27232 5700 27233
rect 5384 27168 5390 27232
rect 5454 27168 5470 27232
rect 5534 27168 5550 27232
rect 5614 27168 5630 27232
rect 5694 27168 5700 27232
rect 5384 27167 5700 27168
rect 9823 27232 10139 27233
rect 9823 27168 9829 27232
rect 9893 27168 9909 27232
rect 9973 27168 9989 27232
rect 10053 27168 10069 27232
rect 10133 27168 10139 27232
rect 9823 27167 10139 27168
rect 14262 27232 14578 27233
rect 14262 27168 14268 27232
rect 14332 27168 14348 27232
rect 14412 27168 14428 27232
rect 14492 27168 14508 27232
rect 14572 27168 14578 27232
rect 14262 27167 14578 27168
rect 18701 27232 19017 27233
rect 18701 27168 18707 27232
rect 18771 27168 18787 27232
rect 18851 27168 18867 27232
rect 18931 27168 18947 27232
rect 19011 27168 19017 27232
rect 18701 27167 19017 27168
rect 7465 27164 7531 27165
rect 7414 27100 7420 27164
rect 7484 27162 7531 27164
rect 7484 27160 7576 27162
rect 7526 27104 7576 27160
rect 7484 27102 7576 27104
rect 7484 27100 7531 27102
rect 7465 27099 7531 27100
rect 0 26754 800 26784
rect 933 26754 999 26757
rect 0 26752 999 26754
rect 0 26696 938 26752
rect 994 26696 999 26752
rect 0 26694 999 26696
rect 0 26664 800 26694
rect 933 26691 999 26694
rect 3165 26688 3481 26689
rect 3165 26624 3171 26688
rect 3235 26624 3251 26688
rect 3315 26624 3331 26688
rect 3395 26624 3411 26688
rect 3475 26624 3481 26688
rect 3165 26623 3481 26624
rect 7604 26688 7920 26689
rect 7604 26624 7610 26688
rect 7674 26624 7690 26688
rect 7754 26624 7770 26688
rect 7834 26624 7850 26688
rect 7914 26624 7920 26688
rect 7604 26623 7920 26624
rect 12043 26688 12359 26689
rect 12043 26624 12049 26688
rect 12113 26624 12129 26688
rect 12193 26624 12209 26688
rect 12273 26624 12289 26688
rect 12353 26624 12359 26688
rect 12043 26623 12359 26624
rect 16482 26688 16798 26689
rect 16482 26624 16488 26688
rect 16552 26624 16568 26688
rect 16632 26624 16648 26688
rect 16712 26624 16728 26688
rect 16792 26624 16798 26688
rect 16482 26623 16798 26624
rect 1761 26618 1827 26621
rect 1894 26618 1900 26620
rect 1761 26616 1900 26618
rect 1761 26560 1766 26616
rect 1822 26560 1900 26616
rect 1761 26558 1900 26560
rect 1761 26555 1827 26558
rect 1894 26556 1900 26558
rect 1964 26556 1970 26620
rect 6177 26346 6243 26349
rect 6678 26346 6684 26348
rect 6177 26344 6684 26346
rect 6177 26288 6182 26344
rect 6238 26288 6684 26344
rect 6177 26286 6684 26288
rect 6177 26283 6243 26286
rect 6678 26284 6684 26286
rect 6748 26284 6754 26348
rect 5384 26144 5700 26145
rect 5384 26080 5390 26144
rect 5454 26080 5470 26144
rect 5534 26080 5550 26144
rect 5614 26080 5630 26144
rect 5694 26080 5700 26144
rect 5384 26079 5700 26080
rect 9823 26144 10139 26145
rect 9823 26080 9829 26144
rect 9893 26080 9909 26144
rect 9973 26080 9989 26144
rect 10053 26080 10069 26144
rect 10133 26080 10139 26144
rect 9823 26079 10139 26080
rect 14262 26144 14578 26145
rect 14262 26080 14268 26144
rect 14332 26080 14348 26144
rect 14412 26080 14428 26144
rect 14492 26080 14508 26144
rect 14572 26080 14578 26144
rect 14262 26079 14578 26080
rect 18701 26144 19017 26145
rect 18701 26080 18707 26144
rect 18771 26080 18787 26144
rect 18851 26080 18867 26144
rect 18931 26080 18947 26144
rect 19011 26080 19017 26144
rect 18701 26079 19017 26080
rect 3165 25600 3481 25601
rect 3165 25536 3171 25600
rect 3235 25536 3251 25600
rect 3315 25536 3331 25600
rect 3395 25536 3411 25600
rect 3475 25536 3481 25600
rect 3165 25535 3481 25536
rect 7604 25600 7920 25601
rect 7604 25536 7610 25600
rect 7674 25536 7690 25600
rect 7754 25536 7770 25600
rect 7834 25536 7850 25600
rect 7914 25536 7920 25600
rect 7604 25535 7920 25536
rect 12043 25600 12359 25601
rect 12043 25536 12049 25600
rect 12113 25536 12129 25600
rect 12193 25536 12209 25600
rect 12273 25536 12289 25600
rect 12353 25536 12359 25600
rect 12043 25535 12359 25536
rect 16482 25600 16798 25601
rect 16482 25536 16488 25600
rect 16552 25536 16568 25600
rect 16632 25536 16648 25600
rect 16712 25536 16728 25600
rect 16792 25536 16798 25600
rect 16482 25535 16798 25536
rect 4838 25196 4844 25260
rect 4908 25258 4914 25260
rect 7833 25258 7899 25261
rect 4908 25256 7899 25258
rect 4908 25200 7838 25256
rect 7894 25200 7899 25256
rect 4908 25198 7899 25200
rect 4908 25196 4914 25198
rect 7833 25195 7899 25198
rect 5384 25056 5700 25057
rect 5384 24992 5390 25056
rect 5454 24992 5470 25056
rect 5534 24992 5550 25056
rect 5614 24992 5630 25056
rect 5694 24992 5700 25056
rect 5384 24991 5700 24992
rect 9823 25056 10139 25057
rect 9823 24992 9829 25056
rect 9893 24992 9909 25056
rect 9973 24992 9989 25056
rect 10053 24992 10069 25056
rect 10133 24992 10139 25056
rect 9823 24991 10139 24992
rect 14262 25056 14578 25057
rect 14262 24992 14268 25056
rect 14332 24992 14348 25056
rect 14412 24992 14428 25056
rect 14492 24992 14508 25056
rect 14572 24992 14578 25056
rect 14262 24991 14578 24992
rect 18701 25056 19017 25057
rect 18701 24992 18707 25056
rect 18771 24992 18787 25056
rect 18851 24992 18867 25056
rect 18931 24992 18947 25056
rect 19011 24992 19017 25056
rect 18701 24991 19017 24992
rect 3165 24512 3481 24513
rect 3165 24448 3171 24512
rect 3235 24448 3251 24512
rect 3315 24448 3331 24512
rect 3395 24448 3411 24512
rect 3475 24448 3481 24512
rect 3165 24447 3481 24448
rect 7604 24512 7920 24513
rect 7604 24448 7610 24512
rect 7674 24448 7690 24512
rect 7754 24448 7770 24512
rect 7834 24448 7850 24512
rect 7914 24448 7920 24512
rect 7604 24447 7920 24448
rect 12043 24512 12359 24513
rect 12043 24448 12049 24512
rect 12113 24448 12129 24512
rect 12193 24448 12209 24512
rect 12273 24448 12289 24512
rect 12353 24448 12359 24512
rect 12043 24447 12359 24448
rect 16482 24512 16798 24513
rect 16482 24448 16488 24512
rect 16552 24448 16568 24512
rect 16632 24448 16648 24512
rect 16712 24448 16728 24512
rect 16792 24448 16798 24512
rect 16482 24447 16798 24448
rect 7005 24170 7071 24173
rect 7414 24170 7420 24172
rect 7005 24168 7420 24170
rect 7005 24112 7010 24168
rect 7066 24112 7420 24168
rect 7005 24110 7420 24112
rect 7005 24107 7071 24110
rect 7414 24108 7420 24110
rect 7484 24108 7490 24172
rect 5384 23968 5700 23969
rect 5384 23904 5390 23968
rect 5454 23904 5470 23968
rect 5534 23904 5550 23968
rect 5614 23904 5630 23968
rect 5694 23904 5700 23968
rect 5384 23903 5700 23904
rect 9823 23968 10139 23969
rect 9823 23904 9829 23968
rect 9893 23904 9909 23968
rect 9973 23904 9989 23968
rect 10053 23904 10069 23968
rect 10133 23904 10139 23968
rect 9823 23903 10139 23904
rect 14262 23968 14578 23969
rect 14262 23904 14268 23968
rect 14332 23904 14348 23968
rect 14412 23904 14428 23968
rect 14492 23904 14508 23968
rect 14572 23904 14578 23968
rect 14262 23903 14578 23904
rect 18701 23968 19017 23969
rect 18701 23904 18707 23968
rect 18771 23904 18787 23968
rect 18851 23904 18867 23968
rect 18931 23904 18947 23968
rect 19011 23904 19017 23968
rect 18701 23903 19017 23904
rect 3918 23428 3924 23492
rect 3988 23490 3994 23492
rect 4061 23490 4127 23493
rect 3988 23488 4127 23490
rect 3988 23432 4066 23488
rect 4122 23432 4127 23488
rect 3988 23430 4127 23432
rect 3988 23428 3994 23430
rect 4061 23427 4127 23430
rect 3165 23424 3481 23425
rect 3165 23360 3171 23424
rect 3235 23360 3251 23424
rect 3315 23360 3331 23424
rect 3395 23360 3411 23424
rect 3475 23360 3481 23424
rect 3165 23359 3481 23360
rect 7604 23424 7920 23425
rect 7604 23360 7610 23424
rect 7674 23360 7690 23424
rect 7754 23360 7770 23424
rect 7834 23360 7850 23424
rect 7914 23360 7920 23424
rect 7604 23359 7920 23360
rect 12043 23424 12359 23425
rect 12043 23360 12049 23424
rect 12113 23360 12129 23424
rect 12193 23360 12209 23424
rect 12273 23360 12289 23424
rect 12353 23360 12359 23424
rect 12043 23359 12359 23360
rect 16482 23424 16798 23425
rect 16482 23360 16488 23424
rect 16552 23360 16568 23424
rect 16632 23360 16648 23424
rect 16712 23360 16728 23424
rect 16792 23360 16798 23424
rect 16482 23359 16798 23360
rect 0 23218 800 23248
rect 933 23218 999 23221
rect 0 23216 999 23218
rect 0 23160 938 23216
rect 994 23160 999 23216
rect 0 23158 999 23160
rect 0 23128 800 23158
rect 933 23155 999 23158
rect 5384 22880 5700 22881
rect 5384 22816 5390 22880
rect 5454 22816 5470 22880
rect 5534 22816 5550 22880
rect 5614 22816 5630 22880
rect 5694 22816 5700 22880
rect 5384 22815 5700 22816
rect 9823 22880 10139 22881
rect 9823 22816 9829 22880
rect 9893 22816 9909 22880
rect 9973 22816 9989 22880
rect 10053 22816 10069 22880
rect 10133 22816 10139 22880
rect 9823 22815 10139 22816
rect 14262 22880 14578 22881
rect 14262 22816 14268 22880
rect 14332 22816 14348 22880
rect 14412 22816 14428 22880
rect 14492 22816 14508 22880
rect 14572 22816 14578 22880
rect 14262 22815 14578 22816
rect 18701 22880 19017 22881
rect 18701 22816 18707 22880
rect 18771 22816 18787 22880
rect 18851 22816 18867 22880
rect 18931 22816 18947 22880
rect 19011 22816 19017 22880
rect 18701 22815 19017 22816
rect 3165 22336 3481 22337
rect 3165 22272 3171 22336
rect 3235 22272 3251 22336
rect 3315 22272 3331 22336
rect 3395 22272 3411 22336
rect 3475 22272 3481 22336
rect 3165 22271 3481 22272
rect 7604 22336 7920 22337
rect 7604 22272 7610 22336
rect 7674 22272 7690 22336
rect 7754 22272 7770 22336
rect 7834 22272 7850 22336
rect 7914 22272 7920 22336
rect 7604 22271 7920 22272
rect 12043 22336 12359 22337
rect 12043 22272 12049 22336
rect 12113 22272 12129 22336
rect 12193 22272 12209 22336
rect 12273 22272 12289 22336
rect 12353 22272 12359 22336
rect 12043 22271 12359 22272
rect 16482 22336 16798 22337
rect 16482 22272 16488 22336
rect 16552 22272 16568 22336
rect 16632 22272 16648 22336
rect 16712 22272 16728 22336
rect 16792 22272 16798 22336
rect 16482 22271 16798 22272
rect 5384 21792 5700 21793
rect 5384 21728 5390 21792
rect 5454 21728 5470 21792
rect 5534 21728 5550 21792
rect 5614 21728 5630 21792
rect 5694 21728 5700 21792
rect 5384 21727 5700 21728
rect 9823 21792 10139 21793
rect 9823 21728 9829 21792
rect 9893 21728 9909 21792
rect 9973 21728 9989 21792
rect 10053 21728 10069 21792
rect 10133 21728 10139 21792
rect 9823 21727 10139 21728
rect 14262 21792 14578 21793
rect 14262 21728 14268 21792
rect 14332 21728 14348 21792
rect 14412 21728 14428 21792
rect 14492 21728 14508 21792
rect 14572 21728 14578 21792
rect 14262 21727 14578 21728
rect 18701 21792 19017 21793
rect 18701 21728 18707 21792
rect 18771 21728 18787 21792
rect 18851 21728 18867 21792
rect 18931 21728 18947 21792
rect 19011 21728 19017 21792
rect 18701 21727 19017 21728
rect 3165 21248 3481 21249
rect 3165 21184 3171 21248
rect 3235 21184 3251 21248
rect 3315 21184 3331 21248
rect 3395 21184 3411 21248
rect 3475 21184 3481 21248
rect 3165 21183 3481 21184
rect 7604 21248 7920 21249
rect 7604 21184 7610 21248
rect 7674 21184 7690 21248
rect 7754 21184 7770 21248
rect 7834 21184 7850 21248
rect 7914 21184 7920 21248
rect 7604 21183 7920 21184
rect 12043 21248 12359 21249
rect 12043 21184 12049 21248
rect 12113 21184 12129 21248
rect 12193 21184 12209 21248
rect 12273 21184 12289 21248
rect 12353 21184 12359 21248
rect 12043 21183 12359 21184
rect 16482 21248 16798 21249
rect 16482 21184 16488 21248
rect 16552 21184 16568 21248
rect 16632 21184 16648 21248
rect 16712 21184 16728 21248
rect 16792 21184 16798 21248
rect 16482 21183 16798 21184
rect 6821 20770 6887 20773
rect 8150 20770 8156 20772
rect 6821 20768 8156 20770
rect 6821 20712 6826 20768
rect 6882 20712 8156 20768
rect 6821 20710 8156 20712
rect 6821 20707 6887 20710
rect 8150 20708 8156 20710
rect 8220 20708 8226 20772
rect 5384 20704 5700 20705
rect 5384 20640 5390 20704
rect 5454 20640 5470 20704
rect 5534 20640 5550 20704
rect 5614 20640 5630 20704
rect 5694 20640 5700 20704
rect 5384 20639 5700 20640
rect 9823 20704 10139 20705
rect 9823 20640 9829 20704
rect 9893 20640 9909 20704
rect 9973 20640 9989 20704
rect 10053 20640 10069 20704
rect 10133 20640 10139 20704
rect 9823 20639 10139 20640
rect 14262 20704 14578 20705
rect 14262 20640 14268 20704
rect 14332 20640 14348 20704
rect 14412 20640 14428 20704
rect 14492 20640 14508 20704
rect 14572 20640 14578 20704
rect 14262 20639 14578 20640
rect 18701 20704 19017 20705
rect 18701 20640 18707 20704
rect 18771 20640 18787 20704
rect 18851 20640 18867 20704
rect 18931 20640 18947 20704
rect 19011 20640 19017 20704
rect 18701 20639 19017 20640
rect 3165 20160 3481 20161
rect 3165 20096 3171 20160
rect 3235 20096 3251 20160
rect 3315 20096 3331 20160
rect 3395 20096 3411 20160
rect 3475 20096 3481 20160
rect 3165 20095 3481 20096
rect 7604 20160 7920 20161
rect 7604 20096 7610 20160
rect 7674 20096 7690 20160
rect 7754 20096 7770 20160
rect 7834 20096 7850 20160
rect 7914 20096 7920 20160
rect 7604 20095 7920 20096
rect 12043 20160 12359 20161
rect 12043 20096 12049 20160
rect 12113 20096 12129 20160
rect 12193 20096 12209 20160
rect 12273 20096 12289 20160
rect 12353 20096 12359 20160
rect 12043 20095 12359 20096
rect 16482 20160 16798 20161
rect 16482 20096 16488 20160
rect 16552 20096 16568 20160
rect 16632 20096 16648 20160
rect 16712 20096 16728 20160
rect 16792 20096 16798 20160
rect 16482 20095 16798 20096
rect 0 19682 800 19712
rect 933 19682 999 19685
rect 0 19680 999 19682
rect 0 19624 938 19680
rect 994 19624 999 19680
rect 0 19622 999 19624
rect 0 19592 800 19622
rect 933 19619 999 19622
rect 5384 19616 5700 19617
rect 5384 19552 5390 19616
rect 5454 19552 5470 19616
rect 5534 19552 5550 19616
rect 5614 19552 5630 19616
rect 5694 19552 5700 19616
rect 5384 19551 5700 19552
rect 9823 19616 10139 19617
rect 9823 19552 9829 19616
rect 9893 19552 9909 19616
rect 9973 19552 9989 19616
rect 10053 19552 10069 19616
rect 10133 19552 10139 19616
rect 9823 19551 10139 19552
rect 14262 19616 14578 19617
rect 14262 19552 14268 19616
rect 14332 19552 14348 19616
rect 14412 19552 14428 19616
rect 14492 19552 14508 19616
rect 14572 19552 14578 19616
rect 14262 19551 14578 19552
rect 18701 19616 19017 19617
rect 18701 19552 18707 19616
rect 18771 19552 18787 19616
rect 18851 19552 18867 19616
rect 18931 19552 18947 19616
rect 19011 19552 19017 19616
rect 18701 19551 19017 19552
rect 2037 19412 2103 19413
rect 2037 19408 2084 19412
rect 2148 19410 2154 19412
rect 2037 19352 2042 19408
rect 2037 19348 2084 19352
rect 2148 19350 2194 19410
rect 2148 19348 2154 19350
rect 2037 19347 2103 19348
rect 3165 19072 3481 19073
rect 3165 19008 3171 19072
rect 3235 19008 3251 19072
rect 3315 19008 3331 19072
rect 3395 19008 3411 19072
rect 3475 19008 3481 19072
rect 3165 19007 3481 19008
rect 7604 19072 7920 19073
rect 7604 19008 7610 19072
rect 7674 19008 7690 19072
rect 7754 19008 7770 19072
rect 7834 19008 7850 19072
rect 7914 19008 7920 19072
rect 7604 19007 7920 19008
rect 12043 19072 12359 19073
rect 12043 19008 12049 19072
rect 12113 19008 12129 19072
rect 12193 19008 12209 19072
rect 12273 19008 12289 19072
rect 12353 19008 12359 19072
rect 12043 19007 12359 19008
rect 16482 19072 16798 19073
rect 16482 19008 16488 19072
rect 16552 19008 16568 19072
rect 16632 19008 16648 19072
rect 16712 19008 16728 19072
rect 16792 19008 16798 19072
rect 16482 19007 16798 19008
rect 5384 18528 5700 18529
rect 5384 18464 5390 18528
rect 5454 18464 5470 18528
rect 5534 18464 5550 18528
rect 5614 18464 5630 18528
rect 5694 18464 5700 18528
rect 5384 18463 5700 18464
rect 9823 18528 10139 18529
rect 9823 18464 9829 18528
rect 9893 18464 9909 18528
rect 9973 18464 9989 18528
rect 10053 18464 10069 18528
rect 10133 18464 10139 18528
rect 9823 18463 10139 18464
rect 14262 18528 14578 18529
rect 14262 18464 14268 18528
rect 14332 18464 14348 18528
rect 14412 18464 14428 18528
rect 14492 18464 14508 18528
rect 14572 18464 14578 18528
rect 14262 18463 14578 18464
rect 18701 18528 19017 18529
rect 18701 18464 18707 18528
rect 18771 18464 18787 18528
rect 18851 18464 18867 18528
rect 18931 18464 18947 18528
rect 19011 18464 19017 18528
rect 18701 18463 19017 18464
rect 3165 17984 3481 17985
rect 3165 17920 3171 17984
rect 3235 17920 3251 17984
rect 3315 17920 3331 17984
rect 3395 17920 3411 17984
rect 3475 17920 3481 17984
rect 3165 17919 3481 17920
rect 7604 17984 7920 17985
rect 7604 17920 7610 17984
rect 7674 17920 7690 17984
rect 7754 17920 7770 17984
rect 7834 17920 7850 17984
rect 7914 17920 7920 17984
rect 7604 17919 7920 17920
rect 12043 17984 12359 17985
rect 12043 17920 12049 17984
rect 12113 17920 12129 17984
rect 12193 17920 12209 17984
rect 12273 17920 12289 17984
rect 12353 17920 12359 17984
rect 12043 17919 12359 17920
rect 16482 17984 16798 17985
rect 16482 17920 16488 17984
rect 16552 17920 16568 17984
rect 16632 17920 16648 17984
rect 16712 17920 16728 17984
rect 16792 17920 16798 17984
rect 16482 17919 16798 17920
rect 5384 17440 5700 17441
rect 5384 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5700 17440
rect 5384 17375 5700 17376
rect 9823 17440 10139 17441
rect 9823 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10139 17440
rect 9823 17375 10139 17376
rect 14262 17440 14578 17441
rect 14262 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14578 17440
rect 14262 17375 14578 17376
rect 18701 17440 19017 17441
rect 18701 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19017 17440
rect 18701 17375 19017 17376
rect 3969 17236 4035 17237
rect 3918 17172 3924 17236
rect 3988 17234 4035 17236
rect 3988 17232 4080 17234
rect 4030 17176 4080 17232
rect 3988 17174 4080 17176
rect 3988 17172 4035 17174
rect 3969 17171 4035 17172
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 16482 16831 16798 16832
rect 2998 16628 3004 16692
rect 3068 16690 3074 16692
rect 3141 16690 3207 16693
rect 3068 16688 3207 16690
rect 3068 16632 3146 16688
rect 3202 16632 3207 16688
rect 3068 16630 3207 16632
rect 3068 16628 3074 16630
rect 3141 16627 3207 16630
rect 5384 16352 5700 16353
rect 5384 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5700 16352
rect 5384 16287 5700 16288
rect 9823 16352 10139 16353
rect 9823 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10139 16352
rect 9823 16287 10139 16288
rect 14262 16352 14578 16353
rect 14262 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14578 16352
rect 14262 16287 14578 16288
rect 18701 16352 19017 16353
rect 18701 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19017 16352
rect 18701 16287 19017 16288
rect 0 16146 800 16176
rect 933 16146 999 16149
rect 0 16144 999 16146
rect 0 16088 938 16144
rect 994 16088 999 16144
rect 0 16086 999 16088
rect 0 16056 800 16086
rect 933 16083 999 16086
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 5384 15264 5700 15265
rect 5384 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5700 15264
rect 5384 15199 5700 15200
rect 9823 15264 10139 15265
rect 9823 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10139 15264
rect 9823 15199 10139 15200
rect 14262 15264 14578 15265
rect 14262 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14578 15264
rect 14262 15199 14578 15200
rect 18701 15264 19017 15265
rect 18701 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19017 15264
rect 18701 15199 19017 15200
rect 3165 14720 3481 14721
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 5384 14176 5700 14177
rect 5384 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5700 14176
rect 5384 14111 5700 14112
rect 9823 14176 10139 14177
rect 9823 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10139 14176
rect 9823 14111 10139 14112
rect 14262 14176 14578 14177
rect 14262 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14578 14176
rect 14262 14111 14578 14112
rect 18701 14176 19017 14177
rect 18701 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19017 14176
rect 18701 14111 19017 14112
rect 2078 13772 2084 13836
rect 2148 13834 2154 13836
rect 5165 13834 5231 13837
rect 2148 13832 5231 13834
rect 2148 13776 5170 13832
rect 5226 13776 5231 13832
rect 2148 13774 5231 13776
rect 2148 13772 2154 13774
rect 5165 13771 5231 13774
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 16482 13567 16798 13568
rect 5384 13088 5700 13089
rect 5384 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5700 13088
rect 5384 13023 5700 13024
rect 9823 13088 10139 13089
rect 9823 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10139 13088
rect 9823 13023 10139 13024
rect 14262 13088 14578 13089
rect 14262 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14578 13088
rect 14262 13023 14578 13024
rect 18701 13088 19017 13089
rect 18701 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19017 13088
rect 18701 13023 19017 13024
rect 3601 12882 3667 12885
rect 3558 12880 3667 12882
rect 3558 12824 3606 12880
rect 3662 12824 3667 12880
rect 3558 12819 3667 12824
rect 2773 12746 2839 12749
rect 3558 12746 3618 12819
rect 2773 12744 3618 12746
rect 2773 12688 2778 12744
rect 2834 12688 3618 12744
rect 2773 12686 3618 12688
rect 2773 12683 2839 12686
rect 0 12610 800 12640
rect 933 12610 999 12613
rect 0 12608 999 12610
rect 0 12552 938 12608
rect 994 12552 999 12608
rect 0 12550 999 12552
rect 0 12520 800 12550
rect 933 12547 999 12550
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 5384 12000 5700 12001
rect 5384 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5700 12000
rect 5384 11935 5700 11936
rect 9823 12000 10139 12001
rect 9823 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10139 12000
rect 9823 11935 10139 11936
rect 14262 12000 14578 12001
rect 14262 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14578 12000
rect 14262 11935 14578 11936
rect 18701 12000 19017 12001
rect 18701 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19017 12000
rect 18701 11935 19017 11936
rect 1894 11596 1900 11660
rect 1964 11658 1970 11660
rect 3601 11658 3667 11661
rect 1964 11656 3667 11658
rect 1964 11600 3606 11656
rect 3662 11600 3667 11656
rect 1964 11598 3667 11600
rect 1964 11596 1970 11598
rect 3601 11595 3667 11598
rect 3165 11456 3481 11457
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 4245 10980 4311 10981
rect 4245 10976 4292 10980
rect 4356 10978 4362 10980
rect 4245 10920 4250 10976
rect 4245 10916 4292 10920
rect 4356 10918 4402 10978
rect 4356 10916 4362 10918
rect 4245 10915 4311 10916
rect 5384 10912 5700 10913
rect 5384 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5700 10912
rect 5384 10847 5700 10848
rect 9823 10912 10139 10913
rect 9823 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10139 10912
rect 9823 10847 10139 10848
rect 14262 10912 14578 10913
rect 14262 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14578 10912
rect 14262 10847 14578 10848
rect 18701 10912 19017 10913
rect 18701 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19017 10912
rect 18701 10847 19017 10848
rect 3165 10368 3481 10369
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 16482 10303 16798 10304
rect 5384 9824 5700 9825
rect 5384 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5700 9824
rect 5384 9759 5700 9760
rect 9823 9824 10139 9825
rect 9823 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10139 9824
rect 9823 9759 10139 9760
rect 14262 9824 14578 9825
rect 14262 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14578 9824
rect 14262 9759 14578 9760
rect 18701 9824 19017 9825
rect 18701 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19017 9824
rect 18701 9759 19017 9760
rect 2773 9754 2839 9757
rect 2998 9754 3004 9756
rect 2773 9752 3004 9754
rect 2773 9696 2778 9752
rect 2834 9696 3004 9752
rect 2773 9694 3004 9696
rect 2773 9691 2839 9694
rect 2998 9692 3004 9694
rect 3068 9692 3074 9756
rect 4061 9618 4127 9621
rect 4654 9618 4660 9620
rect 4061 9616 4660 9618
rect 4061 9560 4066 9616
rect 4122 9560 4660 9616
rect 4061 9558 4660 9560
rect 4061 9555 4127 9558
rect 4654 9556 4660 9558
rect 4724 9556 4730 9620
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 16482 9215 16798 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 5384 8736 5700 8737
rect 5384 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5700 8736
rect 5384 8671 5700 8672
rect 9823 8736 10139 8737
rect 9823 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10139 8736
rect 9823 8671 10139 8672
rect 14262 8736 14578 8737
rect 14262 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14578 8736
rect 14262 8671 14578 8672
rect 18701 8736 19017 8737
rect 18701 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19017 8736
rect 18701 8671 19017 8672
rect 3165 8192 3481 8193
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 2681 6762 2747 6765
rect 2638 6760 2747 6762
rect 2638 6704 2686 6760
rect 2742 6704 2747 6760
rect 2638 6699 2747 6704
rect 2638 6493 2698 6699
rect 6678 6564 6684 6628
rect 6748 6626 6754 6628
rect 6821 6626 6887 6629
rect 6748 6624 6887 6626
rect 6748 6568 6826 6624
rect 6882 6568 6887 6624
rect 6748 6566 6887 6568
rect 6748 6564 6754 6566
rect 6821 6563 6887 6566
rect 5384 6560 5700 6561
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 2589 6488 2698 6493
rect 2589 6432 2594 6488
rect 2650 6432 2698 6488
rect 2589 6430 2698 6432
rect 2589 6427 2655 6430
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 4797 5540 4863 5541
rect 4797 5536 4844 5540
rect 4908 5538 4914 5540
rect 4797 5480 4802 5536
rect 4797 5476 4844 5480
rect 4908 5478 4954 5538
rect 4908 5476 4914 5478
rect 4797 5475 4863 5476
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 18701 5407 19017 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 5384 3296 5700 3297
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 18701 2143 19017 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
<< via3 >>
rect 3171 47356 3235 47360
rect 3171 47300 3175 47356
rect 3175 47300 3231 47356
rect 3231 47300 3235 47356
rect 3171 47296 3235 47300
rect 3251 47356 3315 47360
rect 3251 47300 3255 47356
rect 3255 47300 3311 47356
rect 3311 47300 3315 47356
rect 3251 47296 3315 47300
rect 3331 47356 3395 47360
rect 3331 47300 3335 47356
rect 3335 47300 3391 47356
rect 3391 47300 3395 47356
rect 3331 47296 3395 47300
rect 3411 47356 3475 47360
rect 3411 47300 3415 47356
rect 3415 47300 3471 47356
rect 3471 47300 3475 47356
rect 3411 47296 3475 47300
rect 7610 47356 7674 47360
rect 7610 47300 7614 47356
rect 7614 47300 7670 47356
rect 7670 47300 7674 47356
rect 7610 47296 7674 47300
rect 7690 47356 7754 47360
rect 7690 47300 7694 47356
rect 7694 47300 7750 47356
rect 7750 47300 7754 47356
rect 7690 47296 7754 47300
rect 7770 47356 7834 47360
rect 7770 47300 7774 47356
rect 7774 47300 7830 47356
rect 7830 47300 7834 47356
rect 7770 47296 7834 47300
rect 7850 47356 7914 47360
rect 7850 47300 7854 47356
rect 7854 47300 7910 47356
rect 7910 47300 7914 47356
rect 7850 47296 7914 47300
rect 12049 47356 12113 47360
rect 12049 47300 12053 47356
rect 12053 47300 12109 47356
rect 12109 47300 12113 47356
rect 12049 47296 12113 47300
rect 12129 47356 12193 47360
rect 12129 47300 12133 47356
rect 12133 47300 12189 47356
rect 12189 47300 12193 47356
rect 12129 47296 12193 47300
rect 12209 47356 12273 47360
rect 12209 47300 12213 47356
rect 12213 47300 12269 47356
rect 12269 47300 12273 47356
rect 12209 47296 12273 47300
rect 12289 47356 12353 47360
rect 12289 47300 12293 47356
rect 12293 47300 12349 47356
rect 12349 47300 12353 47356
rect 12289 47296 12353 47300
rect 16488 47356 16552 47360
rect 16488 47300 16492 47356
rect 16492 47300 16548 47356
rect 16548 47300 16552 47356
rect 16488 47296 16552 47300
rect 16568 47356 16632 47360
rect 16568 47300 16572 47356
rect 16572 47300 16628 47356
rect 16628 47300 16632 47356
rect 16568 47296 16632 47300
rect 16648 47356 16712 47360
rect 16648 47300 16652 47356
rect 16652 47300 16708 47356
rect 16708 47300 16712 47356
rect 16648 47296 16712 47300
rect 16728 47356 16792 47360
rect 16728 47300 16732 47356
rect 16732 47300 16788 47356
rect 16788 47300 16792 47356
rect 16728 47296 16792 47300
rect 5390 46812 5454 46816
rect 5390 46756 5394 46812
rect 5394 46756 5450 46812
rect 5450 46756 5454 46812
rect 5390 46752 5454 46756
rect 5470 46812 5534 46816
rect 5470 46756 5474 46812
rect 5474 46756 5530 46812
rect 5530 46756 5534 46812
rect 5470 46752 5534 46756
rect 5550 46812 5614 46816
rect 5550 46756 5554 46812
rect 5554 46756 5610 46812
rect 5610 46756 5614 46812
rect 5550 46752 5614 46756
rect 5630 46812 5694 46816
rect 5630 46756 5634 46812
rect 5634 46756 5690 46812
rect 5690 46756 5694 46812
rect 5630 46752 5694 46756
rect 9829 46812 9893 46816
rect 9829 46756 9833 46812
rect 9833 46756 9889 46812
rect 9889 46756 9893 46812
rect 9829 46752 9893 46756
rect 9909 46812 9973 46816
rect 9909 46756 9913 46812
rect 9913 46756 9969 46812
rect 9969 46756 9973 46812
rect 9909 46752 9973 46756
rect 9989 46812 10053 46816
rect 9989 46756 9993 46812
rect 9993 46756 10049 46812
rect 10049 46756 10053 46812
rect 9989 46752 10053 46756
rect 10069 46812 10133 46816
rect 10069 46756 10073 46812
rect 10073 46756 10129 46812
rect 10129 46756 10133 46812
rect 10069 46752 10133 46756
rect 14268 46812 14332 46816
rect 14268 46756 14272 46812
rect 14272 46756 14328 46812
rect 14328 46756 14332 46812
rect 14268 46752 14332 46756
rect 14348 46812 14412 46816
rect 14348 46756 14352 46812
rect 14352 46756 14408 46812
rect 14408 46756 14412 46812
rect 14348 46752 14412 46756
rect 14428 46812 14492 46816
rect 14428 46756 14432 46812
rect 14432 46756 14488 46812
rect 14488 46756 14492 46812
rect 14428 46752 14492 46756
rect 14508 46812 14572 46816
rect 14508 46756 14512 46812
rect 14512 46756 14568 46812
rect 14568 46756 14572 46812
rect 14508 46752 14572 46756
rect 18707 46812 18771 46816
rect 18707 46756 18711 46812
rect 18711 46756 18767 46812
rect 18767 46756 18771 46812
rect 18707 46752 18771 46756
rect 18787 46812 18851 46816
rect 18787 46756 18791 46812
rect 18791 46756 18847 46812
rect 18847 46756 18851 46812
rect 18787 46752 18851 46756
rect 18867 46812 18931 46816
rect 18867 46756 18871 46812
rect 18871 46756 18927 46812
rect 18927 46756 18931 46812
rect 18867 46752 18931 46756
rect 18947 46812 19011 46816
rect 18947 46756 18951 46812
rect 18951 46756 19007 46812
rect 19007 46756 19011 46812
rect 18947 46752 19011 46756
rect 3171 46268 3235 46272
rect 3171 46212 3175 46268
rect 3175 46212 3231 46268
rect 3231 46212 3235 46268
rect 3171 46208 3235 46212
rect 3251 46268 3315 46272
rect 3251 46212 3255 46268
rect 3255 46212 3311 46268
rect 3311 46212 3315 46268
rect 3251 46208 3315 46212
rect 3331 46268 3395 46272
rect 3331 46212 3335 46268
rect 3335 46212 3391 46268
rect 3391 46212 3395 46268
rect 3331 46208 3395 46212
rect 3411 46268 3475 46272
rect 3411 46212 3415 46268
rect 3415 46212 3471 46268
rect 3471 46212 3475 46268
rect 3411 46208 3475 46212
rect 7610 46268 7674 46272
rect 7610 46212 7614 46268
rect 7614 46212 7670 46268
rect 7670 46212 7674 46268
rect 7610 46208 7674 46212
rect 7690 46268 7754 46272
rect 7690 46212 7694 46268
rect 7694 46212 7750 46268
rect 7750 46212 7754 46268
rect 7690 46208 7754 46212
rect 7770 46268 7834 46272
rect 7770 46212 7774 46268
rect 7774 46212 7830 46268
rect 7830 46212 7834 46268
rect 7770 46208 7834 46212
rect 7850 46268 7914 46272
rect 7850 46212 7854 46268
rect 7854 46212 7910 46268
rect 7910 46212 7914 46268
rect 7850 46208 7914 46212
rect 12049 46268 12113 46272
rect 12049 46212 12053 46268
rect 12053 46212 12109 46268
rect 12109 46212 12113 46268
rect 12049 46208 12113 46212
rect 12129 46268 12193 46272
rect 12129 46212 12133 46268
rect 12133 46212 12189 46268
rect 12189 46212 12193 46268
rect 12129 46208 12193 46212
rect 12209 46268 12273 46272
rect 12209 46212 12213 46268
rect 12213 46212 12269 46268
rect 12269 46212 12273 46268
rect 12209 46208 12273 46212
rect 12289 46268 12353 46272
rect 12289 46212 12293 46268
rect 12293 46212 12349 46268
rect 12349 46212 12353 46268
rect 12289 46208 12353 46212
rect 16488 46268 16552 46272
rect 16488 46212 16492 46268
rect 16492 46212 16548 46268
rect 16548 46212 16552 46268
rect 16488 46208 16552 46212
rect 16568 46268 16632 46272
rect 16568 46212 16572 46268
rect 16572 46212 16628 46268
rect 16628 46212 16632 46268
rect 16568 46208 16632 46212
rect 16648 46268 16712 46272
rect 16648 46212 16652 46268
rect 16652 46212 16708 46268
rect 16708 46212 16712 46268
rect 16648 46208 16712 46212
rect 16728 46268 16792 46272
rect 16728 46212 16732 46268
rect 16732 46212 16788 46268
rect 16788 46212 16792 46268
rect 16728 46208 16792 46212
rect 5390 45724 5454 45728
rect 5390 45668 5394 45724
rect 5394 45668 5450 45724
rect 5450 45668 5454 45724
rect 5390 45664 5454 45668
rect 5470 45724 5534 45728
rect 5470 45668 5474 45724
rect 5474 45668 5530 45724
rect 5530 45668 5534 45724
rect 5470 45664 5534 45668
rect 5550 45724 5614 45728
rect 5550 45668 5554 45724
rect 5554 45668 5610 45724
rect 5610 45668 5614 45724
rect 5550 45664 5614 45668
rect 5630 45724 5694 45728
rect 5630 45668 5634 45724
rect 5634 45668 5690 45724
rect 5690 45668 5694 45724
rect 5630 45664 5694 45668
rect 9829 45724 9893 45728
rect 9829 45668 9833 45724
rect 9833 45668 9889 45724
rect 9889 45668 9893 45724
rect 9829 45664 9893 45668
rect 9909 45724 9973 45728
rect 9909 45668 9913 45724
rect 9913 45668 9969 45724
rect 9969 45668 9973 45724
rect 9909 45664 9973 45668
rect 9989 45724 10053 45728
rect 9989 45668 9993 45724
rect 9993 45668 10049 45724
rect 10049 45668 10053 45724
rect 9989 45664 10053 45668
rect 10069 45724 10133 45728
rect 10069 45668 10073 45724
rect 10073 45668 10129 45724
rect 10129 45668 10133 45724
rect 10069 45664 10133 45668
rect 14268 45724 14332 45728
rect 14268 45668 14272 45724
rect 14272 45668 14328 45724
rect 14328 45668 14332 45724
rect 14268 45664 14332 45668
rect 14348 45724 14412 45728
rect 14348 45668 14352 45724
rect 14352 45668 14408 45724
rect 14408 45668 14412 45724
rect 14348 45664 14412 45668
rect 14428 45724 14492 45728
rect 14428 45668 14432 45724
rect 14432 45668 14488 45724
rect 14488 45668 14492 45724
rect 14428 45664 14492 45668
rect 14508 45724 14572 45728
rect 14508 45668 14512 45724
rect 14512 45668 14568 45724
rect 14568 45668 14572 45724
rect 14508 45664 14572 45668
rect 18707 45724 18771 45728
rect 18707 45668 18711 45724
rect 18711 45668 18767 45724
rect 18767 45668 18771 45724
rect 18707 45664 18771 45668
rect 18787 45724 18851 45728
rect 18787 45668 18791 45724
rect 18791 45668 18847 45724
rect 18847 45668 18851 45724
rect 18787 45664 18851 45668
rect 18867 45724 18931 45728
rect 18867 45668 18871 45724
rect 18871 45668 18927 45724
rect 18927 45668 18931 45724
rect 18867 45664 18931 45668
rect 18947 45724 19011 45728
rect 18947 45668 18951 45724
rect 18951 45668 19007 45724
rect 19007 45668 19011 45724
rect 18947 45664 19011 45668
rect 3171 45180 3235 45184
rect 3171 45124 3175 45180
rect 3175 45124 3231 45180
rect 3231 45124 3235 45180
rect 3171 45120 3235 45124
rect 3251 45180 3315 45184
rect 3251 45124 3255 45180
rect 3255 45124 3311 45180
rect 3311 45124 3315 45180
rect 3251 45120 3315 45124
rect 3331 45180 3395 45184
rect 3331 45124 3335 45180
rect 3335 45124 3391 45180
rect 3391 45124 3395 45180
rect 3331 45120 3395 45124
rect 3411 45180 3475 45184
rect 3411 45124 3415 45180
rect 3415 45124 3471 45180
rect 3471 45124 3475 45180
rect 3411 45120 3475 45124
rect 7610 45180 7674 45184
rect 7610 45124 7614 45180
rect 7614 45124 7670 45180
rect 7670 45124 7674 45180
rect 7610 45120 7674 45124
rect 7690 45180 7754 45184
rect 7690 45124 7694 45180
rect 7694 45124 7750 45180
rect 7750 45124 7754 45180
rect 7690 45120 7754 45124
rect 7770 45180 7834 45184
rect 7770 45124 7774 45180
rect 7774 45124 7830 45180
rect 7830 45124 7834 45180
rect 7770 45120 7834 45124
rect 7850 45180 7914 45184
rect 7850 45124 7854 45180
rect 7854 45124 7910 45180
rect 7910 45124 7914 45180
rect 7850 45120 7914 45124
rect 12049 45180 12113 45184
rect 12049 45124 12053 45180
rect 12053 45124 12109 45180
rect 12109 45124 12113 45180
rect 12049 45120 12113 45124
rect 12129 45180 12193 45184
rect 12129 45124 12133 45180
rect 12133 45124 12189 45180
rect 12189 45124 12193 45180
rect 12129 45120 12193 45124
rect 12209 45180 12273 45184
rect 12209 45124 12213 45180
rect 12213 45124 12269 45180
rect 12269 45124 12273 45180
rect 12209 45120 12273 45124
rect 12289 45180 12353 45184
rect 12289 45124 12293 45180
rect 12293 45124 12349 45180
rect 12349 45124 12353 45180
rect 12289 45120 12353 45124
rect 16488 45180 16552 45184
rect 16488 45124 16492 45180
rect 16492 45124 16548 45180
rect 16548 45124 16552 45180
rect 16488 45120 16552 45124
rect 16568 45180 16632 45184
rect 16568 45124 16572 45180
rect 16572 45124 16628 45180
rect 16628 45124 16632 45180
rect 16568 45120 16632 45124
rect 16648 45180 16712 45184
rect 16648 45124 16652 45180
rect 16652 45124 16708 45180
rect 16708 45124 16712 45180
rect 16648 45120 16712 45124
rect 16728 45180 16792 45184
rect 16728 45124 16732 45180
rect 16732 45124 16788 45180
rect 16788 45124 16792 45180
rect 16728 45120 16792 45124
rect 5390 44636 5454 44640
rect 5390 44580 5394 44636
rect 5394 44580 5450 44636
rect 5450 44580 5454 44636
rect 5390 44576 5454 44580
rect 5470 44636 5534 44640
rect 5470 44580 5474 44636
rect 5474 44580 5530 44636
rect 5530 44580 5534 44636
rect 5470 44576 5534 44580
rect 5550 44636 5614 44640
rect 5550 44580 5554 44636
rect 5554 44580 5610 44636
rect 5610 44580 5614 44636
rect 5550 44576 5614 44580
rect 5630 44636 5694 44640
rect 5630 44580 5634 44636
rect 5634 44580 5690 44636
rect 5690 44580 5694 44636
rect 5630 44576 5694 44580
rect 9829 44636 9893 44640
rect 9829 44580 9833 44636
rect 9833 44580 9889 44636
rect 9889 44580 9893 44636
rect 9829 44576 9893 44580
rect 9909 44636 9973 44640
rect 9909 44580 9913 44636
rect 9913 44580 9969 44636
rect 9969 44580 9973 44636
rect 9909 44576 9973 44580
rect 9989 44636 10053 44640
rect 9989 44580 9993 44636
rect 9993 44580 10049 44636
rect 10049 44580 10053 44636
rect 9989 44576 10053 44580
rect 10069 44636 10133 44640
rect 10069 44580 10073 44636
rect 10073 44580 10129 44636
rect 10129 44580 10133 44636
rect 10069 44576 10133 44580
rect 14268 44636 14332 44640
rect 14268 44580 14272 44636
rect 14272 44580 14328 44636
rect 14328 44580 14332 44636
rect 14268 44576 14332 44580
rect 14348 44636 14412 44640
rect 14348 44580 14352 44636
rect 14352 44580 14408 44636
rect 14408 44580 14412 44636
rect 14348 44576 14412 44580
rect 14428 44636 14492 44640
rect 14428 44580 14432 44636
rect 14432 44580 14488 44636
rect 14488 44580 14492 44636
rect 14428 44576 14492 44580
rect 14508 44636 14572 44640
rect 14508 44580 14512 44636
rect 14512 44580 14568 44636
rect 14568 44580 14572 44636
rect 14508 44576 14572 44580
rect 18707 44636 18771 44640
rect 18707 44580 18711 44636
rect 18711 44580 18767 44636
rect 18767 44580 18771 44636
rect 18707 44576 18771 44580
rect 18787 44636 18851 44640
rect 18787 44580 18791 44636
rect 18791 44580 18847 44636
rect 18847 44580 18851 44636
rect 18787 44576 18851 44580
rect 18867 44636 18931 44640
rect 18867 44580 18871 44636
rect 18871 44580 18927 44636
rect 18927 44580 18931 44636
rect 18867 44576 18931 44580
rect 18947 44636 19011 44640
rect 18947 44580 18951 44636
rect 18951 44580 19007 44636
rect 19007 44580 19011 44636
rect 18947 44576 19011 44580
rect 3171 44092 3235 44096
rect 3171 44036 3175 44092
rect 3175 44036 3231 44092
rect 3231 44036 3235 44092
rect 3171 44032 3235 44036
rect 3251 44092 3315 44096
rect 3251 44036 3255 44092
rect 3255 44036 3311 44092
rect 3311 44036 3315 44092
rect 3251 44032 3315 44036
rect 3331 44092 3395 44096
rect 3331 44036 3335 44092
rect 3335 44036 3391 44092
rect 3391 44036 3395 44092
rect 3331 44032 3395 44036
rect 3411 44092 3475 44096
rect 3411 44036 3415 44092
rect 3415 44036 3471 44092
rect 3471 44036 3475 44092
rect 3411 44032 3475 44036
rect 7610 44092 7674 44096
rect 7610 44036 7614 44092
rect 7614 44036 7670 44092
rect 7670 44036 7674 44092
rect 7610 44032 7674 44036
rect 7690 44092 7754 44096
rect 7690 44036 7694 44092
rect 7694 44036 7750 44092
rect 7750 44036 7754 44092
rect 7690 44032 7754 44036
rect 7770 44092 7834 44096
rect 7770 44036 7774 44092
rect 7774 44036 7830 44092
rect 7830 44036 7834 44092
rect 7770 44032 7834 44036
rect 7850 44092 7914 44096
rect 7850 44036 7854 44092
rect 7854 44036 7910 44092
rect 7910 44036 7914 44092
rect 7850 44032 7914 44036
rect 12049 44092 12113 44096
rect 12049 44036 12053 44092
rect 12053 44036 12109 44092
rect 12109 44036 12113 44092
rect 12049 44032 12113 44036
rect 12129 44092 12193 44096
rect 12129 44036 12133 44092
rect 12133 44036 12189 44092
rect 12189 44036 12193 44092
rect 12129 44032 12193 44036
rect 12209 44092 12273 44096
rect 12209 44036 12213 44092
rect 12213 44036 12269 44092
rect 12269 44036 12273 44092
rect 12209 44032 12273 44036
rect 12289 44092 12353 44096
rect 12289 44036 12293 44092
rect 12293 44036 12349 44092
rect 12349 44036 12353 44092
rect 12289 44032 12353 44036
rect 16488 44092 16552 44096
rect 16488 44036 16492 44092
rect 16492 44036 16548 44092
rect 16548 44036 16552 44092
rect 16488 44032 16552 44036
rect 16568 44092 16632 44096
rect 16568 44036 16572 44092
rect 16572 44036 16628 44092
rect 16628 44036 16632 44092
rect 16568 44032 16632 44036
rect 16648 44092 16712 44096
rect 16648 44036 16652 44092
rect 16652 44036 16708 44092
rect 16708 44036 16712 44092
rect 16648 44032 16712 44036
rect 16728 44092 16792 44096
rect 16728 44036 16732 44092
rect 16732 44036 16788 44092
rect 16788 44036 16792 44092
rect 16728 44032 16792 44036
rect 5390 43548 5454 43552
rect 5390 43492 5394 43548
rect 5394 43492 5450 43548
rect 5450 43492 5454 43548
rect 5390 43488 5454 43492
rect 5470 43548 5534 43552
rect 5470 43492 5474 43548
rect 5474 43492 5530 43548
rect 5530 43492 5534 43548
rect 5470 43488 5534 43492
rect 5550 43548 5614 43552
rect 5550 43492 5554 43548
rect 5554 43492 5610 43548
rect 5610 43492 5614 43548
rect 5550 43488 5614 43492
rect 5630 43548 5694 43552
rect 5630 43492 5634 43548
rect 5634 43492 5690 43548
rect 5690 43492 5694 43548
rect 5630 43488 5694 43492
rect 9829 43548 9893 43552
rect 9829 43492 9833 43548
rect 9833 43492 9889 43548
rect 9889 43492 9893 43548
rect 9829 43488 9893 43492
rect 9909 43548 9973 43552
rect 9909 43492 9913 43548
rect 9913 43492 9969 43548
rect 9969 43492 9973 43548
rect 9909 43488 9973 43492
rect 9989 43548 10053 43552
rect 9989 43492 9993 43548
rect 9993 43492 10049 43548
rect 10049 43492 10053 43548
rect 9989 43488 10053 43492
rect 10069 43548 10133 43552
rect 10069 43492 10073 43548
rect 10073 43492 10129 43548
rect 10129 43492 10133 43548
rect 10069 43488 10133 43492
rect 14268 43548 14332 43552
rect 14268 43492 14272 43548
rect 14272 43492 14328 43548
rect 14328 43492 14332 43548
rect 14268 43488 14332 43492
rect 14348 43548 14412 43552
rect 14348 43492 14352 43548
rect 14352 43492 14408 43548
rect 14408 43492 14412 43548
rect 14348 43488 14412 43492
rect 14428 43548 14492 43552
rect 14428 43492 14432 43548
rect 14432 43492 14488 43548
rect 14488 43492 14492 43548
rect 14428 43488 14492 43492
rect 14508 43548 14572 43552
rect 14508 43492 14512 43548
rect 14512 43492 14568 43548
rect 14568 43492 14572 43548
rect 14508 43488 14572 43492
rect 18707 43548 18771 43552
rect 18707 43492 18711 43548
rect 18711 43492 18767 43548
rect 18767 43492 18771 43548
rect 18707 43488 18771 43492
rect 18787 43548 18851 43552
rect 18787 43492 18791 43548
rect 18791 43492 18847 43548
rect 18847 43492 18851 43548
rect 18787 43488 18851 43492
rect 18867 43548 18931 43552
rect 18867 43492 18871 43548
rect 18871 43492 18927 43548
rect 18927 43492 18931 43548
rect 18867 43488 18931 43492
rect 18947 43548 19011 43552
rect 18947 43492 18951 43548
rect 18951 43492 19007 43548
rect 19007 43492 19011 43548
rect 18947 43488 19011 43492
rect 3171 43004 3235 43008
rect 3171 42948 3175 43004
rect 3175 42948 3231 43004
rect 3231 42948 3235 43004
rect 3171 42944 3235 42948
rect 3251 43004 3315 43008
rect 3251 42948 3255 43004
rect 3255 42948 3311 43004
rect 3311 42948 3315 43004
rect 3251 42944 3315 42948
rect 3331 43004 3395 43008
rect 3331 42948 3335 43004
rect 3335 42948 3391 43004
rect 3391 42948 3395 43004
rect 3331 42944 3395 42948
rect 3411 43004 3475 43008
rect 3411 42948 3415 43004
rect 3415 42948 3471 43004
rect 3471 42948 3475 43004
rect 3411 42944 3475 42948
rect 7610 43004 7674 43008
rect 7610 42948 7614 43004
rect 7614 42948 7670 43004
rect 7670 42948 7674 43004
rect 7610 42944 7674 42948
rect 7690 43004 7754 43008
rect 7690 42948 7694 43004
rect 7694 42948 7750 43004
rect 7750 42948 7754 43004
rect 7690 42944 7754 42948
rect 7770 43004 7834 43008
rect 7770 42948 7774 43004
rect 7774 42948 7830 43004
rect 7830 42948 7834 43004
rect 7770 42944 7834 42948
rect 7850 43004 7914 43008
rect 7850 42948 7854 43004
rect 7854 42948 7910 43004
rect 7910 42948 7914 43004
rect 7850 42944 7914 42948
rect 12049 43004 12113 43008
rect 12049 42948 12053 43004
rect 12053 42948 12109 43004
rect 12109 42948 12113 43004
rect 12049 42944 12113 42948
rect 12129 43004 12193 43008
rect 12129 42948 12133 43004
rect 12133 42948 12189 43004
rect 12189 42948 12193 43004
rect 12129 42944 12193 42948
rect 12209 43004 12273 43008
rect 12209 42948 12213 43004
rect 12213 42948 12269 43004
rect 12269 42948 12273 43004
rect 12209 42944 12273 42948
rect 12289 43004 12353 43008
rect 12289 42948 12293 43004
rect 12293 42948 12349 43004
rect 12349 42948 12353 43004
rect 12289 42944 12353 42948
rect 16488 43004 16552 43008
rect 16488 42948 16492 43004
rect 16492 42948 16548 43004
rect 16548 42948 16552 43004
rect 16488 42944 16552 42948
rect 16568 43004 16632 43008
rect 16568 42948 16572 43004
rect 16572 42948 16628 43004
rect 16628 42948 16632 43004
rect 16568 42944 16632 42948
rect 16648 43004 16712 43008
rect 16648 42948 16652 43004
rect 16652 42948 16708 43004
rect 16708 42948 16712 43004
rect 16648 42944 16712 42948
rect 16728 43004 16792 43008
rect 16728 42948 16732 43004
rect 16732 42948 16788 43004
rect 16788 42948 16792 43004
rect 16728 42944 16792 42948
rect 5390 42460 5454 42464
rect 5390 42404 5394 42460
rect 5394 42404 5450 42460
rect 5450 42404 5454 42460
rect 5390 42400 5454 42404
rect 5470 42460 5534 42464
rect 5470 42404 5474 42460
rect 5474 42404 5530 42460
rect 5530 42404 5534 42460
rect 5470 42400 5534 42404
rect 5550 42460 5614 42464
rect 5550 42404 5554 42460
rect 5554 42404 5610 42460
rect 5610 42404 5614 42460
rect 5550 42400 5614 42404
rect 5630 42460 5694 42464
rect 5630 42404 5634 42460
rect 5634 42404 5690 42460
rect 5690 42404 5694 42460
rect 5630 42400 5694 42404
rect 9829 42460 9893 42464
rect 9829 42404 9833 42460
rect 9833 42404 9889 42460
rect 9889 42404 9893 42460
rect 9829 42400 9893 42404
rect 9909 42460 9973 42464
rect 9909 42404 9913 42460
rect 9913 42404 9969 42460
rect 9969 42404 9973 42460
rect 9909 42400 9973 42404
rect 9989 42460 10053 42464
rect 9989 42404 9993 42460
rect 9993 42404 10049 42460
rect 10049 42404 10053 42460
rect 9989 42400 10053 42404
rect 10069 42460 10133 42464
rect 10069 42404 10073 42460
rect 10073 42404 10129 42460
rect 10129 42404 10133 42460
rect 10069 42400 10133 42404
rect 14268 42460 14332 42464
rect 14268 42404 14272 42460
rect 14272 42404 14328 42460
rect 14328 42404 14332 42460
rect 14268 42400 14332 42404
rect 14348 42460 14412 42464
rect 14348 42404 14352 42460
rect 14352 42404 14408 42460
rect 14408 42404 14412 42460
rect 14348 42400 14412 42404
rect 14428 42460 14492 42464
rect 14428 42404 14432 42460
rect 14432 42404 14488 42460
rect 14488 42404 14492 42460
rect 14428 42400 14492 42404
rect 14508 42460 14572 42464
rect 14508 42404 14512 42460
rect 14512 42404 14568 42460
rect 14568 42404 14572 42460
rect 14508 42400 14572 42404
rect 18707 42460 18771 42464
rect 18707 42404 18711 42460
rect 18711 42404 18767 42460
rect 18767 42404 18771 42460
rect 18707 42400 18771 42404
rect 18787 42460 18851 42464
rect 18787 42404 18791 42460
rect 18791 42404 18847 42460
rect 18847 42404 18851 42460
rect 18787 42400 18851 42404
rect 18867 42460 18931 42464
rect 18867 42404 18871 42460
rect 18871 42404 18927 42460
rect 18927 42404 18931 42460
rect 18867 42400 18931 42404
rect 18947 42460 19011 42464
rect 18947 42404 18951 42460
rect 18951 42404 19007 42460
rect 19007 42404 19011 42460
rect 18947 42400 19011 42404
rect 3171 41916 3235 41920
rect 3171 41860 3175 41916
rect 3175 41860 3231 41916
rect 3231 41860 3235 41916
rect 3171 41856 3235 41860
rect 3251 41916 3315 41920
rect 3251 41860 3255 41916
rect 3255 41860 3311 41916
rect 3311 41860 3315 41916
rect 3251 41856 3315 41860
rect 3331 41916 3395 41920
rect 3331 41860 3335 41916
rect 3335 41860 3391 41916
rect 3391 41860 3395 41916
rect 3331 41856 3395 41860
rect 3411 41916 3475 41920
rect 3411 41860 3415 41916
rect 3415 41860 3471 41916
rect 3471 41860 3475 41916
rect 3411 41856 3475 41860
rect 7610 41916 7674 41920
rect 7610 41860 7614 41916
rect 7614 41860 7670 41916
rect 7670 41860 7674 41916
rect 7610 41856 7674 41860
rect 7690 41916 7754 41920
rect 7690 41860 7694 41916
rect 7694 41860 7750 41916
rect 7750 41860 7754 41916
rect 7690 41856 7754 41860
rect 7770 41916 7834 41920
rect 7770 41860 7774 41916
rect 7774 41860 7830 41916
rect 7830 41860 7834 41916
rect 7770 41856 7834 41860
rect 7850 41916 7914 41920
rect 7850 41860 7854 41916
rect 7854 41860 7910 41916
rect 7910 41860 7914 41916
rect 7850 41856 7914 41860
rect 12049 41916 12113 41920
rect 12049 41860 12053 41916
rect 12053 41860 12109 41916
rect 12109 41860 12113 41916
rect 12049 41856 12113 41860
rect 12129 41916 12193 41920
rect 12129 41860 12133 41916
rect 12133 41860 12189 41916
rect 12189 41860 12193 41916
rect 12129 41856 12193 41860
rect 12209 41916 12273 41920
rect 12209 41860 12213 41916
rect 12213 41860 12269 41916
rect 12269 41860 12273 41916
rect 12209 41856 12273 41860
rect 12289 41916 12353 41920
rect 12289 41860 12293 41916
rect 12293 41860 12349 41916
rect 12349 41860 12353 41916
rect 12289 41856 12353 41860
rect 16488 41916 16552 41920
rect 16488 41860 16492 41916
rect 16492 41860 16548 41916
rect 16548 41860 16552 41916
rect 16488 41856 16552 41860
rect 16568 41916 16632 41920
rect 16568 41860 16572 41916
rect 16572 41860 16628 41916
rect 16628 41860 16632 41916
rect 16568 41856 16632 41860
rect 16648 41916 16712 41920
rect 16648 41860 16652 41916
rect 16652 41860 16708 41916
rect 16708 41860 16712 41916
rect 16648 41856 16712 41860
rect 16728 41916 16792 41920
rect 16728 41860 16732 41916
rect 16732 41860 16788 41916
rect 16788 41860 16792 41916
rect 16728 41856 16792 41860
rect 5390 41372 5454 41376
rect 5390 41316 5394 41372
rect 5394 41316 5450 41372
rect 5450 41316 5454 41372
rect 5390 41312 5454 41316
rect 5470 41372 5534 41376
rect 5470 41316 5474 41372
rect 5474 41316 5530 41372
rect 5530 41316 5534 41372
rect 5470 41312 5534 41316
rect 5550 41372 5614 41376
rect 5550 41316 5554 41372
rect 5554 41316 5610 41372
rect 5610 41316 5614 41372
rect 5550 41312 5614 41316
rect 5630 41372 5694 41376
rect 5630 41316 5634 41372
rect 5634 41316 5690 41372
rect 5690 41316 5694 41372
rect 5630 41312 5694 41316
rect 9829 41372 9893 41376
rect 9829 41316 9833 41372
rect 9833 41316 9889 41372
rect 9889 41316 9893 41372
rect 9829 41312 9893 41316
rect 9909 41372 9973 41376
rect 9909 41316 9913 41372
rect 9913 41316 9969 41372
rect 9969 41316 9973 41372
rect 9909 41312 9973 41316
rect 9989 41372 10053 41376
rect 9989 41316 9993 41372
rect 9993 41316 10049 41372
rect 10049 41316 10053 41372
rect 9989 41312 10053 41316
rect 10069 41372 10133 41376
rect 10069 41316 10073 41372
rect 10073 41316 10129 41372
rect 10129 41316 10133 41372
rect 10069 41312 10133 41316
rect 14268 41372 14332 41376
rect 14268 41316 14272 41372
rect 14272 41316 14328 41372
rect 14328 41316 14332 41372
rect 14268 41312 14332 41316
rect 14348 41372 14412 41376
rect 14348 41316 14352 41372
rect 14352 41316 14408 41372
rect 14408 41316 14412 41372
rect 14348 41312 14412 41316
rect 14428 41372 14492 41376
rect 14428 41316 14432 41372
rect 14432 41316 14488 41372
rect 14488 41316 14492 41372
rect 14428 41312 14492 41316
rect 14508 41372 14572 41376
rect 14508 41316 14512 41372
rect 14512 41316 14568 41372
rect 14568 41316 14572 41372
rect 14508 41312 14572 41316
rect 18707 41372 18771 41376
rect 18707 41316 18711 41372
rect 18711 41316 18767 41372
rect 18767 41316 18771 41372
rect 18707 41312 18771 41316
rect 18787 41372 18851 41376
rect 18787 41316 18791 41372
rect 18791 41316 18847 41372
rect 18847 41316 18851 41372
rect 18787 41312 18851 41316
rect 18867 41372 18931 41376
rect 18867 41316 18871 41372
rect 18871 41316 18927 41372
rect 18927 41316 18931 41372
rect 18867 41312 18931 41316
rect 18947 41372 19011 41376
rect 18947 41316 18951 41372
rect 18951 41316 19007 41372
rect 19007 41316 19011 41372
rect 18947 41312 19011 41316
rect 3171 40828 3235 40832
rect 3171 40772 3175 40828
rect 3175 40772 3231 40828
rect 3231 40772 3235 40828
rect 3171 40768 3235 40772
rect 3251 40828 3315 40832
rect 3251 40772 3255 40828
rect 3255 40772 3311 40828
rect 3311 40772 3315 40828
rect 3251 40768 3315 40772
rect 3331 40828 3395 40832
rect 3331 40772 3335 40828
rect 3335 40772 3391 40828
rect 3391 40772 3395 40828
rect 3331 40768 3395 40772
rect 3411 40828 3475 40832
rect 3411 40772 3415 40828
rect 3415 40772 3471 40828
rect 3471 40772 3475 40828
rect 3411 40768 3475 40772
rect 7610 40828 7674 40832
rect 7610 40772 7614 40828
rect 7614 40772 7670 40828
rect 7670 40772 7674 40828
rect 7610 40768 7674 40772
rect 7690 40828 7754 40832
rect 7690 40772 7694 40828
rect 7694 40772 7750 40828
rect 7750 40772 7754 40828
rect 7690 40768 7754 40772
rect 7770 40828 7834 40832
rect 7770 40772 7774 40828
rect 7774 40772 7830 40828
rect 7830 40772 7834 40828
rect 7770 40768 7834 40772
rect 7850 40828 7914 40832
rect 7850 40772 7854 40828
rect 7854 40772 7910 40828
rect 7910 40772 7914 40828
rect 7850 40768 7914 40772
rect 12049 40828 12113 40832
rect 12049 40772 12053 40828
rect 12053 40772 12109 40828
rect 12109 40772 12113 40828
rect 12049 40768 12113 40772
rect 12129 40828 12193 40832
rect 12129 40772 12133 40828
rect 12133 40772 12189 40828
rect 12189 40772 12193 40828
rect 12129 40768 12193 40772
rect 12209 40828 12273 40832
rect 12209 40772 12213 40828
rect 12213 40772 12269 40828
rect 12269 40772 12273 40828
rect 12209 40768 12273 40772
rect 12289 40828 12353 40832
rect 12289 40772 12293 40828
rect 12293 40772 12349 40828
rect 12349 40772 12353 40828
rect 12289 40768 12353 40772
rect 16488 40828 16552 40832
rect 16488 40772 16492 40828
rect 16492 40772 16548 40828
rect 16548 40772 16552 40828
rect 16488 40768 16552 40772
rect 16568 40828 16632 40832
rect 16568 40772 16572 40828
rect 16572 40772 16628 40828
rect 16628 40772 16632 40828
rect 16568 40768 16632 40772
rect 16648 40828 16712 40832
rect 16648 40772 16652 40828
rect 16652 40772 16708 40828
rect 16708 40772 16712 40828
rect 16648 40768 16712 40772
rect 16728 40828 16792 40832
rect 16728 40772 16732 40828
rect 16732 40772 16788 40828
rect 16788 40772 16792 40828
rect 16728 40768 16792 40772
rect 5390 40284 5454 40288
rect 5390 40228 5394 40284
rect 5394 40228 5450 40284
rect 5450 40228 5454 40284
rect 5390 40224 5454 40228
rect 5470 40284 5534 40288
rect 5470 40228 5474 40284
rect 5474 40228 5530 40284
rect 5530 40228 5534 40284
rect 5470 40224 5534 40228
rect 5550 40284 5614 40288
rect 5550 40228 5554 40284
rect 5554 40228 5610 40284
rect 5610 40228 5614 40284
rect 5550 40224 5614 40228
rect 5630 40284 5694 40288
rect 5630 40228 5634 40284
rect 5634 40228 5690 40284
rect 5690 40228 5694 40284
rect 5630 40224 5694 40228
rect 9829 40284 9893 40288
rect 9829 40228 9833 40284
rect 9833 40228 9889 40284
rect 9889 40228 9893 40284
rect 9829 40224 9893 40228
rect 9909 40284 9973 40288
rect 9909 40228 9913 40284
rect 9913 40228 9969 40284
rect 9969 40228 9973 40284
rect 9909 40224 9973 40228
rect 9989 40284 10053 40288
rect 9989 40228 9993 40284
rect 9993 40228 10049 40284
rect 10049 40228 10053 40284
rect 9989 40224 10053 40228
rect 10069 40284 10133 40288
rect 10069 40228 10073 40284
rect 10073 40228 10129 40284
rect 10129 40228 10133 40284
rect 10069 40224 10133 40228
rect 14268 40284 14332 40288
rect 14268 40228 14272 40284
rect 14272 40228 14328 40284
rect 14328 40228 14332 40284
rect 14268 40224 14332 40228
rect 14348 40284 14412 40288
rect 14348 40228 14352 40284
rect 14352 40228 14408 40284
rect 14408 40228 14412 40284
rect 14348 40224 14412 40228
rect 14428 40284 14492 40288
rect 14428 40228 14432 40284
rect 14432 40228 14488 40284
rect 14488 40228 14492 40284
rect 14428 40224 14492 40228
rect 14508 40284 14572 40288
rect 14508 40228 14512 40284
rect 14512 40228 14568 40284
rect 14568 40228 14572 40284
rect 14508 40224 14572 40228
rect 18707 40284 18771 40288
rect 18707 40228 18711 40284
rect 18711 40228 18767 40284
rect 18767 40228 18771 40284
rect 18707 40224 18771 40228
rect 18787 40284 18851 40288
rect 18787 40228 18791 40284
rect 18791 40228 18847 40284
rect 18847 40228 18851 40284
rect 18787 40224 18851 40228
rect 18867 40284 18931 40288
rect 18867 40228 18871 40284
rect 18871 40228 18927 40284
rect 18927 40228 18931 40284
rect 18867 40224 18931 40228
rect 18947 40284 19011 40288
rect 18947 40228 18951 40284
rect 18951 40228 19007 40284
rect 19007 40228 19011 40284
rect 18947 40224 19011 40228
rect 3171 39740 3235 39744
rect 3171 39684 3175 39740
rect 3175 39684 3231 39740
rect 3231 39684 3235 39740
rect 3171 39680 3235 39684
rect 3251 39740 3315 39744
rect 3251 39684 3255 39740
rect 3255 39684 3311 39740
rect 3311 39684 3315 39740
rect 3251 39680 3315 39684
rect 3331 39740 3395 39744
rect 3331 39684 3335 39740
rect 3335 39684 3391 39740
rect 3391 39684 3395 39740
rect 3331 39680 3395 39684
rect 3411 39740 3475 39744
rect 3411 39684 3415 39740
rect 3415 39684 3471 39740
rect 3471 39684 3475 39740
rect 3411 39680 3475 39684
rect 7610 39740 7674 39744
rect 7610 39684 7614 39740
rect 7614 39684 7670 39740
rect 7670 39684 7674 39740
rect 7610 39680 7674 39684
rect 7690 39740 7754 39744
rect 7690 39684 7694 39740
rect 7694 39684 7750 39740
rect 7750 39684 7754 39740
rect 7690 39680 7754 39684
rect 7770 39740 7834 39744
rect 7770 39684 7774 39740
rect 7774 39684 7830 39740
rect 7830 39684 7834 39740
rect 7770 39680 7834 39684
rect 7850 39740 7914 39744
rect 7850 39684 7854 39740
rect 7854 39684 7910 39740
rect 7910 39684 7914 39740
rect 7850 39680 7914 39684
rect 12049 39740 12113 39744
rect 12049 39684 12053 39740
rect 12053 39684 12109 39740
rect 12109 39684 12113 39740
rect 12049 39680 12113 39684
rect 12129 39740 12193 39744
rect 12129 39684 12133 39740
rect 12133 39684 12189 39740
rect 12189 39684 12193 39740
rect 12129 39680 12193 39684
rect 12209 39740 12273 39744
rect 12209 39684 12213 39740
rect 12213 39684 12269 39740
rect 12269 39684 12273 39740
rect 12209 39680 12273 39684
rect 12289 39740 12353 39744
rect 12289 39684 12293 39740
rect 12293 39684 12349 39740
rect 12349 39684 12353 39740
rect 12289 39680 12353 39684
rect 16488 39740 16552 39744
rect 16488 39684 16492 39740
rect 16492 39684 16548 39740
rect 16548 39684 16552 39740
rect 16488 39680 16552 39684
rect 16568 39740 16632 39744
rect 16568 39684 16572 39740
rect 16572 39684 16628 39740
rect 16628 39684 16632 39740
rect 16568 39680 16632 39684
rect 16648 39740 16712 39744
rect 16648 39684 16652 39740
rect 16652 39684 16708 39740
rect 16708 39684 16712 39740
rect 16648 39680 16712 39684
rect 16728 39740 16792 39744
rect 16728 39684 16732 39740
rect 16732 39684 16788 39740
rect 16788 39684 16792 39740
rect 16728 39680 16792 39684
rect 5390 39196 5454 39200
rect 5390 39140 5394 39196
rect 5394 39140 5450 39196
rect 5450 39140 5454 39196
rect 5390 39136 5454 39140
rect 5470 39196 5534 39200
rect 5470 39140 5474 39196
rect 5474 39140 5530 39196
rect 5530 39140 5534 39196
rect 5470 39136 5534 39140
rect 5550 39196 5614 39200
rect 5550 39140 5554 39196
rect 5554 39140 5610 39196
rect 5610 39140 5614 39196
rect 5550 39136 5614 39140
rect 5630 39196 5694 39200
rect 5630 39140 5634 39196
rect 5634 39140 5690 39196
rect 5690 39140 5694 39196
rect 5630 39136 5694 39140
rect 9829 39196 9893 39200
rect 9829 39140 9833 39196
rect 9833 39140 9889 39196
rect 9889 39140 9893 39196
rect 9829 39136 9893 39140
rect 9909 39196 9973 39200
rect 9909 39140 9913 39196
rect 9913 39140 9969 39196
rect 9969 39140 9973 39196
rect 9909 39136 9973 39140
rect 9989 39196 10053 39200
rect 9989 39140 9993 39196
rect 9993 39140 10049 39196
rect 10049 39140 10053 39196
rect 9989 39136 10053 39140
rect 10069 39196 10133 39200
rect 10069 39140 10073 39196
rect 10073 39140 10129 39196
rect 10129 39140 10133 39196
rect 10069 39136 10133 39140
rect 14268 39196 14332 39200
rect 14268 39140 14272 39196
rect 14272 39140 14328 39196
rect 14328 39140 14332 39196
rect 14268 39136 14332 39140
rect 14348 39196 14412 39200
rect 14348 39140 14352 39196
rect 14352 39140 14408 39196
rect 14408 39140 14412 39196
rect 14348 39136 14412 39140
rect 14428 39196 14492 39200
rect 14428 39140 14432 39196
rect 14432 39140 14488 39196
rect 14488 39140 14492 39196
rect 14428 39136 14492 39140
rect 14508 39196 14572 39200
rect 14508 39140 14512 39196
rect 14512 39140 14568 39196
rect 14568 39140 14572 39196
rect 14508 39136 14572 39140
rect 18707 39196 18771 39200
rect 18707 39140 18711 39196
rect 18711 39140 18767 39196
rect 18767 39140 18771 39196
rect 18707 39136 18771 39140
rect 18787 39196 18851 39200
rect 18787 39140 18791 39196
rect 18791 39140 18847 39196
rect 18847 39140 18851 39196
rect 18787 39136 18851 39140
rect 18867 39196 18931 39200
rect 18867 39140 18871 39196
rect 18871 39140 18927 39196
rect 18927 39140 18931 39196
rect 18867 39136 18931 39140
rect 18947 39196 19011 39200
rect 18947 39140 18951 39196
rect 18951 39140 19007 39196
rect 19007 39140 19011 39196
rect 18947 39136 19011 39140
rect 3171 38652 3235 38656
rect 3171 38596 3175 38652
rect 3175 38596 3231 38652
rect 3231 38596 3235 38652
rect 3171 38592 3235 38596
rect 3251 38652 3315 38656
rect 3251 38596 3255 38652
rect 3255 38596 3311 38652
rect 3311 38596 3315 38652
rect 3251 38592 3315 38596
rect 3331 38652 3395 38656
rect 3331 38596 3335 38652
rect 3335 38596 3391 38652
rect 3391 38596 3395 38652
rect 3331 38592 3395 38596
rect 3411 38652 3475 38656
rect 3411 38596 3415 38652
rect 3415 38596 3471 38652
rect 3471 38596 3475 38652
rect 3411 38592 3475 38596
rect 7610 38652 7674 38656
rect 7610 38596 7614 38652
rect 7614 38596 7670 38652
rect 7670 38596 7674 38652
rect 7610 38592 7674 38596
rect 7690 38652 7754 38656
rect 7690 38596 7694 38652
rect 7694 38596 7750 38652
rect 7750 38596 7754 38652
rect 7690 38592 7754 38596
rect 7770 38652 7834 38656
rect 7770 38596 7774 38652
rect 7774 38596 7830 38652
rect 7830 38596 7834 38652
rect 7770 38592 7834 38596
rect 7850 38652 7914 38656
rect 7850 38596 7854 38652
rect 7854 38596 7910 38652
rect 7910 38596 7914 38652
rect 7850 38592 7914 38596
rect 12049 38652 12113 38656
rect 12049 38596 12053 38652
rect 12053 38596 12109 38652
rect 12109 38596 12113 38652
rect 12049 38592 12113 38596
rect 12129 38652 12193 38656
rect 12129 38596 12133 38652
rect 12133 38596 12189 38652
rect 12189 38596 12193 38652
rect 12129 38592 12193 38596
rect 12209 38652 12273 38656
rect 12209 38596 12213 38652
rect 12213 38596 12269 38652
rect 12269 38596 12273 38652
rect 12209 38592 12273 38596
rect 12289 38652 12353 38656
rect 12289 38596 12293 38652
rect 12293 38596 12349 38652
rect 12349 38596 12353 38652
rect 12289 38592 12353 38596
rect 16488 38652 16552 38656
rect 16488 38596 16492 38652
rect 16492 38596 16548 38652
rect 16548 38596 16552 38652
rect 16488 38592 16552 38596
rect 16568 38652 16632 38656
rect 16568 38596 16572 38652
rect 16572 38596 16628 38652
rect 16628 38596 16632 38652
rect 16568 38592 16632 38596
rect 16648 38652 16712 38656
rect 16648 38596 16652 38652
rect 16652 38596 16708 38652
rect 16708 38596 16712 38652
rect 16648 38592 16712 38596
rect 16728 38652 16792 38656
rect 16728 38596 16732 38652
rect 16732 38596 16788 38652
rect 16788 38596 16792 38652
rect 16728 38592 16792 38596
rect 5390 38108 5454 38112
rect 5390 38052 5394 38108
rect 5394 38052 5450 38108
rect 5450 38052 5454 38108
rect 5390 38048 5454 38052
rect 5470 38108 5534 38112
rect 5470 38052 5474 38108
rect 5474 38052 5530 38108
rect 5530 38052 5534 38108
rect 5470 38048 5534 38052
rect 5550 38108 5614 38112
rect 5550 38052 5554 38108
rect 5554 38052 5610 38108
rect 5610 38052 5614 38108
rect 5550 38048 5614 38052
rect 5630 38108 5694 38112
rect 5630 38052 5634 38108
rect 5634 38052 5690 38108
rect 5690 38052 5694 38108
rect 5630 38048 5694 38052
rect 9829 38108 9893 38112
rect 9829 38052 9833 38108
rect 9833 38052 9889 38108
rect 9889 38052 9893 38108
rect 9829 38048 9893 38052
rect 9909 38108 9973 38112
rect 9909 38052 9913 38108
rect 9913 38052 9969 38108
rect 9969 38052 9973 38108
rect 9909 38048 9973 38052
rect 9989 38108 10053 38112
rect 9989 38052 9993 38108
rect 9993 38052 10049 38108
rect 10049 38052 10053 38108
rect 9989 38048 10053 38052
rect 10069 38108 10133 38112
rect 10069 38052 10073 38108
rect 10073 38052 10129 38108
rect 10129 38052 10133 38108
rect 10069 38048 10133 38052
rect 14268 38108 14332 38112
rect 14268 38052 14272 38108
rect 14272 38052 14328 38108
rect 14328 38052 14332 38108
rect 14268 38048 14332 38052
rect 14348 38108 14412 38112
rect 14348 38052 14352 38108
rect 14352 38052 14408 38108
rect 14408 38052 14412 38108
rect 14348 38048 14412 38052
rect 14428 38108 14492 38112
rect 14428 38052 14432 38108
rect 14432 38052 14488 38108
rect 14488 38052 14492 38108
rect 14428 38048 14492 38052
rect 14508 38108 14572 38112
rect 14508 38052 14512 38108
rect 14512 38052 14568 38108
rect 14568 38052 14572 38108
rect 14508 38048 14572 38052
rect 18707 38108 18771 38112
rect 18707 38052 18711 38108
rect 18711 38052 18767 38108
rect 18767 38052 18771 38108
rect 18707 38048 18771 38052
rect 18787 38108 18851 38112
rect 18787 38052 18791 38108
rect 18791 38052 18847 38108
rect 18847 38052 18851 38108
rect 18787 38048 18851 38052
rect 18867 38108 18931 38112
rect 18867 38052 18871 38108
rect 18871 38052 18927 38108
rect 18927 38052 18931 38108
rect 18867 38048 18931 38052
rect 18947 38108 19011 38112
rect 18947 38052 18951 38108
rect 18951 38052 19007 38108
rect 19007 38052 19011 38108
rect 18947 38048 19011 38052
rect 3171 37564 3235 37568
rect 3171 37508 3175 37564
rect 3175 37508 3231 37564
rect 3231 37508 3235 37564
rect 3171 37504 3235 37508
rect 3251 37564 3315 37568
rect 3251 37508 3255 37564
rect 3255 37508 3311 37564
rect 3311 37508 3315 37564
rect 3251 37504 3315 37508
rect 3331 37564 3395 37568
rect 3331 37508 3335 37564
rect 3335 37508 3391 37564
rect 3391 37508 3395 37564
rect 3331 37504 3395 37508
rect 3411 37564 3475 37568
rect 3411 37508 3415 37564
rect 3415 37508 3471 37564
rect 3471 37508 3475 37564
rect 3411 37504 3475 37508
rect 7610 37564 7674 37568
rect 7610 37508 7614 37564
rect 7614 37508 7670 37564
rect 7670 37508 7674 37564
rect 7610 37504 7674 37508
rect 7690 37564 7754 37568
rect 7690 37508 7694 37564
rect 7694 37508 7750 37564
rect 7750 37508 7754 37564
rect 7690 37504 7754 37508
rect 7770 37564 7834 37568
rect 7770 37508 7774 37564
rect 7774 37508 7830 37564
rect 7830 37508 7834 37564
rect 7770 37504 7834 37508
rect 7850 37564 7914 37568
rect 7850 37508 7854 37564
rect 7854 37508 7910 37564
rect 7910 37508 7914 37564
rect 7850 37504 7914 37508
rect 12049 37564 12113 37568
rect 12049 37508 12053 37564
rect 12053 37508 12109 37564
rect 12109 37508 12113 37564
rect 12049 37504 12113 37508
rect 12129 37564 12193 37568
rect 12129 37508 12133 37564
rect 12133 37508 12189 37564
rect 12189 37508 12193 37564
rect 12129 37504 12193 37508
rect 12209 37564 12273 37568
rect 12209 37508 12213 37564
rect 12213 37508 12269 37564
rect 12269 37508 12273 37564
rect 12209 37504 12273 37508
rect 12289 37564 12353 37568
rect 12289 37508 12293 37564
rect 12293 37508 12349 37564
rect 12349 37508 12353 37564
rect 12289 37504 12353 37508
rect 16488 37564 16552 37568
rect 16488 37508 16492 37564
rect 16492 37508 16548 37564
rect 16548 37508 16552 37564
rect 16488 37504 16552 37508
rect 16568 37564 16632 37568
rect 16568 37508 16572 37564
rect 16572 37508 16628 37564
rect 16628 37508 16632 37564
rect 16568 37504 16632 37508
rect 16648 37564 16712 37568
rect 16648 37508 16652 37564
rect 16652 37508 16708 37564
rect 16708 37508 16712 37564
rect 16648 37504 16712 37508
rect 16728 37564 16792 37568
rect 16728 37508 16732 37564
rect 16732 37508 16788 37564
rect 16788 37508 16792 37564
rect 16728 37504 16792 37508
rect 5390 37020 5454 37024
rect 5390 36964 5394 37020
rect 5394 36964 5450 37020
rect 5450 36964 5454 37020
rect 5390 36960 5454 36964
rect 5470 37020 5534 37024
rect 5470 36964 5474 37020
rect 5474 36964 5530 37020
rect 5530 36964 5534 37020
rect 5470 36960 5534 36964
rect 5550 37020 5614 37024
rect 5550 36964 5554 37020
rect 5554 36964 5610 37020
rect 5610 36964 5614 37020
rect 5550 36960 5614 36964
rect 5630 37020 5694 37024
rect 5630 36964 5634 37020
rect 5634 36964 5690 37020
rect 5690 36964 5694 37020
rect 5630 36960 5694 36964
rect 9829 37020 9893 37024
rect 9829 36964 9833 37020
rect 9833 36964 9889 37020
rect 9889 36964 9893 37020
rect 9829 36960 9893 36964
rect 9909 37020 9973 37024
rect 9909 36964 9913 37020
rect 9913 36964 9969 37020
rect 9969 36964 9973 37020
rect 9909 36960 9973 36964
rect 9989 37020 10053 37024
rect 9989 36964 9993 37020
rect 9993 36964 10049 37020
rect 10049 36964 10053 37020
rect 9989 36960 10053 36964
rect 10069 37020 10133 37024
rect 10069 36964 10073 37020
rect 10073 36964 10129 37020
rect 10129 36964 10133 37020
rect 10069 36960 10133 36964
rect 14268 37020 14332 37024
rect 14268 36964 14272 37020
rect 14272 36964 14328 37020
rect 14328 36964 14332 37020
rect 14268 36960 14332 36964
rect 14348 37020 14412 37024
rect 14348 36964 14352 37020
rect 14352 36964 14408 37020
rect 14408 36964 14412 37020
rect 14348 36960 14412 36964
rect 14428 37020 14492 37024
rect 14428 36964 14432 37020
rect 14432 36964 14488 37020
rect 14488 36964 14492 37020
rect 14428 36960 14492 36964
rect 14508 37020 14572 37024
rect 14508 36964 14512 37020
rect 14512 36964 14568 37020
rect 14568 36964 14572 37020
rect 14508 36960 14572 36964
rect 18707 37020 18771 37024
rect 18707 36964 18711 37020
rect 18711 36964 18767 37020
rect 18767 36964 18771 37020
rect 18707 36960 18771 36964
rect 18787 37020 18851 37024
rect 18787 36964 18791 37020
rect 18791 36964 18847 37020
rect 18847 36964 18851 37020
rect 18787 36960 18851 36964
rect 18867 37020 18931 37024
rect 18867 36964 18871 37020
rect 18871 36964 18927 37020
rect 18927 36964 18931 37020
rect 18867 36960 18931 36964
rect 18947 37020 19011 37024
rect 18947 36964 18951 37020
rect 18951 36964 19007 37020
rect 19007 36964 19011 37020
rect 18947 36960 19011 36964
rect 3171 36476 3235 36480
rect 3171 36420 3175 36476
rect 3175 36420 3231 36476
rect 3231 36420 3235 36476
rect 3171 36416 3235 36420
rect 3251 36476 3315 36480
rect 3251 36420 3255 36476
rect 3255 36420 3311 36476
rect 3311 36420 3315 36476
rect 3251 36416 3315 36420
rect 3331 36476 3395 36480
rect 3331 36420 3335 36476
rect 3335 36420 3391 36476
rect 3391 36420 3395 36476
rect 3331 36416 3395 36420
rect 3411 36476 3475 36480
rect 3411 36420 3415 36476
rect 3415 36420 3471 36476
rect 3471 36420 3475 36476
rect 3411 36416 3475 36420
rect 7610 36476 7674 36480
rect 7610 36420 7614 36476
rect 7614 36420 7670 36476
rect 7670 36420 7674 36476
rect 7610 36416 7674 36420
rect 7690 36476 7754 36480
rect 7690 36420 7694 36476
rect 7694 36420 7750 36476
rect 7750 36420 7754 36476
rect 7690 36416 7754 36420
rect 7770 36476 7834 36480
rect 7770 36420 7774 36476
rect 7774 36420 7830 36476
rect 7830 36420 7834 36476
rect 7770 36416 7834 36420
rect 7850 36476 7914 36480
rect 7850 36420 7854 36476
rect 7854 36420 7910 36476
rect 7910 36420 7914 36476
rect 7850 36416 7914 36420
rect 12049 36476 12113 36480
rect 12049 36420 12053 36476
rect 12053 36420 12109 36476
rect 12109 36420 12113 36476
rect 12049 36416 12113 36420
rect 12129 36476 12193 36480
rect 12129 36420 12133 36476
rect 12133 36420 12189 36476
rect 12189 36420 12193 36476
rect 12129 36416 12193 36420
rect 12209 36476 12273 36480
rect 12209 36420 12213 36476
rect 12213 36420 12269 36476
rect 12269 36420 12273 36476
rect 12209 36416 12273 36420
rect 12289 36476 12353 36480
rect 12289 36420 12293 36476
rect 12293 36420 12349 36476
rect 12349 36420 12353 36476
rect 12289 36416 12353 36420
rect 16488 36476 16552 36480
rect 16488 36420 16492 36476
rect 16492 36420 16548 36476
rect 16548 36420 16552 36476
rect 16488 36416 16552 36420
rect 16568 36476 16632 36480
rect 16568 36420 16572 36476
rect 16572 36420 16628 36476
rect 16628 36420 16632 36476
rect 16568 36416 16632 36420
rect 16648 36476 16712 36480
rect 16648 36420 16652 36476
rect 16652 36420 16708 36476
rect 16708 36420 16712 36476
rect 16648 36416 16712 36420
rect 16728 36476 16792 36480
rect 16728 36420 16732 36476
rect 16732 36420 16788 36476
rect 16788 36420 16792 36476
rect 16728 36416 16792 36420
rect 5390 35932 5454 35936
rect 5390 35876 5394 35932
rect 5394 35876 5450 35932
rect 5450 35876 5454 35932
rect 5390 35872 5454 35876
rect 5470 35932 5534 35936
rect 5470 35876 5474 35932
rect 5474 35876 5530 35932
rect 5530 35876 5534 35932
rect 5470 35872 5534 35876
rect 5550 35932 5614 35936
rect 5550 35876 5554 35932
rect 5554 35876 5610 35932
rect 5610 35876 5614 35932
rect 5550 35872 5614 35876
rect 5630 35932 5694 35936
rect 5630 35876 5634 35932
rect 5634 35876 5690 35932
rect 5690 35876 5694 35932
rect 5630 35872 5694 35876
rect 9829 35932 9893 35936
rect 9829 35876 9833 35932
rect 9833 35876 9889 35932
rect 9889 35876 9893 35932
rect 9829 35872 9893 35876
rect 9909 35932 9973 35936
rect 9909 35876 9913 35932
rect 9913 35876 9969 35932
rect 9969 35876 9973 35932
rect 9909 35872 9973 35876
rect 9989 35932 10053 35936
rect 9989 35876 9993 35932
rect 9993 35876 10049 35932
rect 10049 35876 10053 35932
rect 9989 35872 10053 35876
rect 10069 35932 10133 35936
rect 10069 35876 10073 35932
rect 10073 35876 10129 35932
rect 10129 35876 10133 35932
rect 10069 35872 10133 35876
rect 14268 35932 14332 35936
rect 14268 35876 14272 35932
rect 14272 35876 14328 35932
rect 14328 35876 14332 35932
rect 14268 35872 14332 35876
rect 14348 35932 14412 35936
rect 14348 35876 14352 35932
rect 14352 35876 14408 35932
rect 14408 35876 14412 35932
rect 14348 35872 14412 35876
rect 14428 35932 14492 35936
rect 14428 35876 14432 35932
rect 14432 35876 14488 35932
rect 14488 35876 14492 35932
rect 14428 35872 14492 35876
rect 14508 35932 14572 35936
rect 14508 35876 14512 35932
rect 14512 35876 14568 35932
rect 14568 35876 14572 35932
rect 14508 35872 14572 35876
rect 18707 35932 18771 35936
rect 18707 35876 18711 35932
rect 18711 35876 18767 35932
rect 18767 35876 18771 35932
rect 18707 35872 18771 35876
rect 18787 35932 18851 35936
rect 18787 35876 18791 35932
rect 18791 35876 18847 35932
rect 18847 35876 18851 35932
rect 18787 35872 18851 35876
rect 18867 35932 18931 35936
rect 18867 35876 18871 35932
rect 18871 35876 18927 35932
rect 18927 35876 18931 35932
rect 18867 35872 18931 35876
rect 18947 35932 19011 35936
rect 18947 35876 18951 35932
rect 18951 35876 19007 35932
rect 19007 35876 19011 35932
rect 18947 35872 19011 35876
rect 3171 35388 3235 35392
rect 3171 35332 3175 35388
rect 3175 35332 3231 35388
rect 3231 35332 3235 35388
rect 3171 35328 3235 35332
rect 3251 35388 3315 35392
rect 3251 35332 3255 35388
rect 3255 35332 3311 35388
rect 3311 35332 3315 35388
rect 3251 35328 3315 35332
rect 3331 35388 3395 35392
rect 3331 35332 3335 35388
rect 3335 35332 3391 35388
rect 3391 35332 3395 35388
rect 3331 35328 3395 35332
rect 3411 35388 3475 35392
rect 3411 35332 3415 35388
rect 3415 35332 3471 35388
rect 3471 35332 3475 35388
rect 3411 35328 3475 35332
rect 7610 35388 7674 35392
rect 7610 35332 7614 35388
rect 7614 35332 7670 35388
rect 7670 35332 7674 35388
rect 7610 35328 7674 35332
rect 7690 35388 7754 35392
rect 7690 35332 7694 35388
rect 7694 35332 7750 35388
rect 7750 35332 7754 35388
rect 7690 35328 7754 35332
rect 7770 35388 7834 35392
rect 7770 35332 7774 35388
rect 7774 35332 7830 35388
rect 7830 35332 7834 35388
rect 7770 35328 7834 35332
rect 7850 35388 7914 35392
rect 7850 35332 7854 35388
rect 7854 35332 7910 35388
rect 7910 35332 7914 35388
rect 7850 35328 7914 35332
rect 12049 35388 12113 35392
rect 12049 35332 12053 35388
rect 12053 35332 12109 35388
rect 12109 35332 12113 35388
rect 12049 35328 12113 35332
rect 12129 35388 12193 35392
rect 12129 35332 12133 35388
rect 12133 35332 12189 35388
rect 12189 35332 12193 35388
rect 12129 35328 12193 35332
rect 12209 35388 12273 35392
rect 12209 35332 12213 35388
rect 12213 35332 12269 35388
rect 12269 35332 12273 35388
rect 12209 35328 12273 35332
rect 12289 35388 12353 35392
rect 12289 35332 12293 35388
rect 12293 35332 12349 35388
rect 12349 35332 12353 35388
rect 12289 35328 12353 35332
rect 16488 35388 16552 35392
rect 16488 35332 16492 35388
rect 16492 35332 16548 35388
rect 16548 35332 16552 35388
rect 16488 35328 16552 35332
rect 16568 35388 16632 35392
rect 16568 35332 16572 35388
rect 16572 35332 16628 35388
rect 16628 35332 16632 35388
rect 16568 35328 16632 35332
rect 16648 35388 16712 35392
rect 16648 35332 16652 35388
rect 16652 35332 16708 35388
rect 16708 35332 16712 35388
rect 16648 35328 16712 35332
rect 16728 35388 16792 35392
rect 16728 35332 16732 35388
rect 16732 35332 16788 35388
rect 16788 35332 16792 35388
rect 16728 35328 16792 35332
rect 5390 34844 5454 34848
rect 5390 34788 5394 34844
rect 5394 34788 5450 34844
rect 5450 34788 5454 34844
rect 5390 34784 5454 34788
rect 5470 34844 5534 34848
rect 5470 34788 5474 34844
rect 5474 34788 5530 34844
rect 5530 34788 5534 34844
rect 5470 34784 5534 34788
rect 5550 34844 5614 34848
rect 5550 34788 5554 34844
rect 5554 34788 5610 34844
rect 5610 34788 5614 34844
rect 5550 34784 5614 34788
rect 5630 34844 5694 34848
rect 5630 34788 5634 34844
rect 5634 34788 5690 34844
rect 5690 34788 5694 34844
rect 5630 34784 5694 34788
rect 9829 34844 9893 34848
rect 9829 34788 9833 34844
rect 9833 34788 9889 34844
rect 9889 34788 9893 34844
rect 9829 34784 9893 34788
rect 9909 34844 9973 34848
rect 9909 34788 9913 34844
rect 9913 34788 9969 34844
rect 9969 34788 9973 34844
rect 9909 34784 9973 34788
rect 9989 34844 10053 34848
rect 9989 34788 9993 34844
rect 9993 34788 10049 34844
rect 10049 34788 10053 34844
rect 9989 34784 10053 34788
rect 10069 34844 10133 34848
rect 10069 34788 10073 34844
rect 10073 34788 10129 34844
rect 10129 34788 10133 34844
rect 10069 34784 10133 34788
rect 14268 34844 14332 34848
rect 14268 34788 14272 34844
rect 14272 34788 14328 34844
rect 14328 34788 14332 34844
rect 14268 34784 14332 34788
rect 14348 34844 14412 34848
rect 14348 34788 14352 34844
rect 14352 34788 14408 34844
rect 14408 34788 14412 34844
rect 14348 34784 14412 34788
rect 14428 34844 14492 34848
rect 14428 34788 14432 34844
rect 14432 34788 14488 34844
rect 14488 34788 14492 34844
rect 14428 34784 14492 34788
rect 14508 34844 14572 34848
rect 14508 34788 14512 34844
rect 14512 34788 14568 34844
rect 14568 34788 14572 34844
rect 14508 34784 14572 34788
rect 18707 34844 18771 34848
rect 18707 34788 18711 34844
rect 18711 34788 18767 34844
rect 18767 34788 18771 34844
rect 18707 34784 18771 34788
rect 18787 34844 18851 34848
rect 18787 34788 18791 34844
rect 18791 34788 18847 34844
rect 18847 34788 18851 34844
rect 18787 34784 18851 34788
rect 18867 34844 18931 34848
rect 18867 34788 18871 34844
rect 18871 34788 18927 34844
rect 18927 34788 18931 34844
rect 18867 34784 18931 34788
rect 18947 34844 19011 34848
rect 18947 34788 18951 34844
rect 18951 34788 19007 34844
rect 19007 34788 19011 34844
rect 18947 34784 19011 34788
rect 3171 34300 3235 34304
rect 3171 34244 3175 34300
rect 3175 34244 3231 34300
rect 3231 34244 3235 34300
rect 3171 34240 3235 34244
rect 3251 34300 3315 34304
rect 3251 34244 3255 34300
rect 3255 34244 3311 34300
rect 3311 34244 3315 34300
rect 3251 34240 3315 34244
rect 3331 34300 3395 34304
rect 3331 34244 3335 34300
rect 3335 34244 3391 34300
rect 3391 34244 3395 34300
rect 3331 34240 3395 34244
rect 3411 34300 3475 34304
rect 3411 34244 3415 34300
rect 3415 34244 3471 34300
rect 3471 34244 3475 34300
rect 3411 34240 3475 34244
rect 7610 34300 7674 34304
rect 7610 34244 7614 34300
rect 7614 34244 7670 34300
rect 7670 34244 7674 34300
rect 7610 34240 7674 34244
rect 7690 34300 7754 34304
rect 7690 34244 7694 34300
rect 7694 34244 7750 34300
rect 7750 34244 7754 34300
rect 7690 34240 7754 34244
rect 7770 34300 7834 34304
rect 7770 34244 7774 34300
rect 7774 34244 7830 34300
rect 7830 34244 7834 34300
rect 7770 34240 7834 34244
rect 7850 34300 7914 34304
rect 7850 34244 7854 34300
rect 7854 34244 7910 34300
rect 7910 34244 7914 34300
rect 7850 34240 7914 34244
rect 12049 34300 12113 34304
rect 12049 34244 12053 34300
rect 12053 34244 12109 34300
rect 12109 34244 12113 34300
rect 12049 34240 12113 34244
rect 12129 34300 12193 34304
rect 12129 34244 12133 34300
rect 12133 34244 12189 34300
rect 12189 34244 12193 34300
rect 12129 34240 12193 34244
rect 12209 34300 12273 34304
rect 12209 34244 12213 34300
rect 12213 34244 12269 34300
rect 12269 34244 12273 34300
rect 12209 34240 12273 34244
rect 12289 34300 12353 34304
rect 12289 34244 12293 34300
rect 12293 34244 12349 34300
rect 12349 34244 12353 34300
rect 12289 34240 12353 34244
rect 16488 34300 16552 34304
rect 16488 34244 16492 34300
rect 16492 34244 16548 34300
rect 16548 34244 16552 34300
rect 16488 34240 16552 34244
rect 16568 34300 16632 34304
rect 16568 34244 16572 34300
rect 16572 34244 16628 34300
rect 16628 34244 16632 34300
rect 16568 34240 16632 34244
rect 16648 34300 16712 34304
rect 16648 34244 16652 34300
rect 16652 34244 16708 34300
rect 16708 34244 16712 34300
rect 16648 34240 16712 34244
rect 16728 34300 16792 34304
rect 16728 34244 16732 34300
rect 16732 34244 16788 34300
rect 16788 34244 16792 34300
rect 16728 34240 16792 34244
rect 5390 33756 5454 33760
rect 5390 33700 5394 33756
rect 5394 33700 5450 33756
rect 5450 33700 5454 33756
rect 5390 33696 5454 33700
rect 5470 33756 5534 33760
rect 5470 33700 5474 33756
rect 5474 33700 5530 33756
rect 5530 33700 5534 33756
rect 5470 33696 5534 33700
rect 5550 33756 5614 33760
rect 5550 33700 5554 33756
rect 5554 33700 5610 33756
rect 5610 33700 5614 33756
rect 5550 33696 5614 33700
rect 5630 33756 5694 33760
rect 5630 33700 5634 33756
rect 5634 33700 5690 33756
rect 5690 33700 5694 33756
rect 5630 33696 5694 33700
rect 9829 33756 9893 33760
rect 9829 33700 9833 33756
rect 9833 33700 9889 33756
rect 9889 33700 9893 33756
rect 9829 33696 9893 33700
rect 9909 33756 9973 33760
rect 9909 33700 9913 33756
rect 9913 33700 9969 33756
rect 9969 33700 9973 33756
rect 9909 33696 9973 33700
rect 9989 33756 10053 33760
rect 9989 33700 9993 33756
rect 9993 33700 10049 33756
rect 10049 33700 10053 33756
rect 9989 33696 10053 33700
rect 10069 33756 10133 33760
rect 10069 33700 10073 33756
rect 10073 33700 10129 33756
rect 10129 33700 10133 33756
rect 10069 33696 10133 33700
rect 14268 33756 14332 33760
rect 14268 33700 14272 33756
rect 14272 33700 14328 33756
rect 14328 33700 14332 33756
rect 14268 33696 14332 33700
rect 14348 33756 14412 33760
rect 14348 33700 14352 33756
rect 14352 33700 14408 33756
rect 14408 33700 14412 33756
rect 14348 33696 14412 33700
rect 14428 33756 14492 33760
rect 14428 33700 14432 33756
rect 14432 33700 14488 33756
rect 14488 33700 14492 33756
rect 14428 33696 14492 33700
rect 14508 33756 14572 33760
rect 14508 33700 14512 33756
rect 14512 33700 14568 33756
rect 14568 33700 14572 33756
rect 14508 33696 14572 33700
rect 18707 33756 18771 33760
rect 18707 33700 18711 33756
rect 18711 33700 18767 33756
rect 18767 33700 18771 33756
rect 18707 33696 18771 33700
rect 18787 33756 18851 33760
rect 18787 33700 18791 33756
rect 18791 33700 18847 33756
rect 18847 33700 18851 33756
rect 18787 33696 18851 33700
rect 18867 33756 18931 33760
rect 18867 33700 18871 33756
rect 18871 33700 18927 33756
rect 18927 33700 18931 33756
rect 18867 33696 18931 33700
rect 18947 33756 19011 33760
rect 18947 33700 18951 33756
rect 18951 33700 19007 33756
rect 19007 33700 19011 33756
rect 18947 33696 19011 33700
rect 3171 33212 3235 33216
rect 3171 33156 3175 33212
rect 3175 33156 3231 33212
rect 3231 33156 3235 33212
rect 3171 33152 3235 33156
rect 3251 33212 3315 33216
rect 3251 33156 3255 33212
rect 3255 33156 3311 33212
rect 3311 33156 3315 33212
rect 3251 33152 3315 33156
rect 3331 33212 3395 33216
rect 3331 33156 3335 33212
rect 3335 33156 3391 33212
rect 3391 33156 3395 33212
rect 3331 33152 3395 33156
rect 3411 33212 3475 33216
rect 3411 33156 3415 33212
rect 3415 33156 3471 33212
rect 3471 33156 3475 33212
rect 3411 33152 3475 33156
rect 7610 33212 7674 33216
rect 7610 33156 7614 33212
rect 7614 33156 7670 33212
rect 7670 33156 7674 33212
rect 7610 33152 7674 33156
rect 7690 33212 7754 33216
rect 7690 33156 7694 33212
rect 7694 33156 7750 33212
rect 7750 33156 7754 33212
rect 7690 33152 7754 33156
rect 7770 33212 7834 33216
rect 7770 33156 7774 33212
rect 7774 33156 7830 33212
rect 7830 33156 7834 33212
rect 7770 33152 7834 33156
rect 7850 33212 7914 33216
rect 7850 33156 7854 33212
rect 7854 33156 7910 33212
rect 7910 33156 7914 33212
rect 7850 33152 7914 33156
rect 12049 33212 12113 33216
rect 12049 33156 12053 33212
rect 12053 33156 12109 33212
rect 12109 33156 12113 33212
rect 12049 33152 12113 33156
rect 12129 33212 12193 33216
rect 12129 33156 12133 33212
rect 12133 33156 12189 33212
rect 12189 33156 12193 33212
rect 12129 33152 12193 33156
rect 12209 33212 12273 33216
rect 12209 33156 12213 33212
rect 12213 33156 12269 33212
rect 12269 33156 12273 33212
rect 12209 33152 12273 33156
rect 12289 33212 12353 33216
rect 12289 33156 12293 33212
rect 12293 33156 12349 33212
rect 12349 33156 12353 33212
rect 12289 33152 12353 33156
rect 16488 33212 16552 33216
rect 16488 33156 16492 33212
rect 16492 33156 16548 33212
rect 16548 33156 16552 33212
rect 16488 33152 16552 33156
rect 16568 33212 16632 33216
rect 16568 33156 16572 33212
rect 16572 33156 16628 33212
rect 16628 33156 16632 33212
rect 16568 33152 16632 33156
rect 16648 33212 16712 33216
rect 16648 33156 16652 33212
rect 16652 33156 16708 33212
rect 16708 33156 16712 33212
rect 16648 33152 16712 33156
rect 16728 33212 16792 33216
rect 16728 33156 16732 33212
rect 16732 33156 16788 33212
rect 16788 33156 16792 33212
rect 16728 33152 16792 33156
rect 5390 32668 5454 32672
rect 5390 32612 5394 32668
rect 5394 32612 5450 32668
rect 5450 32612 5454 32668
rect 5390 32608 5454 32612
rect 5470 32668 5534 32672
rect 5470 32612 5474 32668
rect 5474 32612 5530 32668
rect 5530 32612 5534 32668
rect 5470 32608 5534 32612
rect 5550 32668 5614 32672
rect 5550 32612 5554 32668
rect 5554 32612 5610 32668
rect 5610 32612 5614 32668
rect 5550 32608 5614 32612
rect 5630 32668 5694 32672
rect 5630 32612 5634 32668
rect 5634 32612 5690 32668
rect 5690 32612 5694 32668
rect 5630 32608 5694 32612
rect 9829 32668 9893 32672
rect 9829 32612 9833 32668
rect 9833 32612 9889 32668
rect 9889 32612 9893 32668
rect 9829 32608 9893 32612
rect 9909 32668 9973 32672
rect 9909 32612 9913 32668
rect 9913 32612 9969 32668
rect 9969 32612 9973 32668
rect 9909 32608 9973 32612
rect 9989 32668 10053 32672
rect 9989 32612 9993 32668
rect 9993 32612 10049 32668
rect 10049 32612 10053 32668
rect 9989 32608 10053 32612
rect 10069 32668 10133 32672
rect 10069 32612 10073 32668
rect 10073 32612 10129 32668
rect 10129 32612 10133 32668
rect 10069 32608 10133 32612
rect 14268 32668 14332 32672
rect 14268 32612 14272 32668
rect 14272 32612 14328 32668
rect 14328 32612 14332 32668
rect 14268 32608 14332 32612
rect 14348 32668 14412 32672
rect 14348 32612 14352 32668
rect 14352 32612 14408 32668
rect 14408 32612 14412 32668
rect 14348 32608 14412 32612
rect 14428 32668 14492 32672
rect 14428 32612 14432 32668
rect 14432 32612 14488 32668
rect 14488 32612 14492 32668
rect 14428 32608 14492 32612
rect 14508 32668 14572 32672
rect 14508 32612 14512 32668
rect 14512 32612 14568 32668
rect 14568 32612 14572 32668
rect 14508 32608 14572 32612
rect 18707 32668 18771 32672
rect 18707 32612 18711 32668
rect 18711 32612 18767 32668
rect 18767 32612 18771 32668
rect 18707 32608 18771 32612
rect 18787 32668 18851 32672
rect 18787 32612 18791 32668
rect 18791 32612 18847 32668
rect 18847 32612 18851 32668
rect 18787 32608 18851 32612
rect 18867 32668 18931 32672
rect 18867 32612 18871 32668
rect 18871 32612 18927 32668
rect 18927 32612 18931 32668
rect 18867 32608 18931 32612
rect 18947 32668 19011 32672
rect 18947 32612 18951 32668
rect 18951 32612 19007 32668
rect 19007 32612 19011 32668
rect 18947 32608 19011 32612
rect 3171 32124 3235 32128
rect 3171 32068 3175 32124
rect 3175 32068 3231 32124
rect 3231 32068 3235 32124
rect 3171 32064 3235 32068
rect 3251 32124 3315 32128
rect 3251 32068 3255 32124
rect 3255 32068 3311 32124
rect 3311 32068 3315 32124
rect 3251 32064 3315 32068
rect 3331 32124 3395 32128
rect 3331 32068 3335 32124
rect 3335 32068 3391 32124
rect 3391 32068 3395 32124
rect 3331 32064 3395 32068
rect 3411 32124 3475 32128
rect 3411 32068 3415 32124
rect 3415 32068 3471 32124
rect 3471 32068 3475 32124
rect 3411 32064 3475 32068
rect 7610 32124 7674 32128
rect 7610 32068 7614 32124
rect 7614 32068 7670 32124
rect 7670 32068 7674 32124
rect 7610 32064 7674 32068
rect 7690 32124 7754 32128
rect 7690 32068 7694 32124
rect 7694 32068 7750 32124
rect 7750 32068 7754 32124
rect 7690 32064 7754 32068
rect 7770 32124 7834 32128
rect 7770 32068 7774 32124
rect 7774 32068 7830 32124
rect 7830 32068 7834 32124
rect 7770 32064 7834 32068
rect 7850 32124 7914 32128
rect 7850 32068 7854 32124
rect 7854 32068 7910 32124
rect 7910 32068 7914 32124
rect 7850 32064 7914 32068
rect 12049 32124 12113 32128
rect 12049 32068 12053 32124
rect 12053 32068 12109 32124
rect 12109 32068 12113 32124
rect 12049 32064 12113 32068
rect 12129 32124 12193 32128
rect 12129 32068 12133 32124
rect 12133 32068 12189 32124
rect 12189 32068 12193 32124
rect 12129 32064 12193 32068
rect 12209 32124 12273 32128
rect 12209 32068 12213 32124
rect 12213 32068 12269 32124
rect 12269 32068 12273 32124
rect 12209 32064 12273 32068
rect 12289 32124 12353 32128
rect 12289 32068 12293 32124
rect 12293 32068 12349 32124
rect 12349 32068 12353 32124
rect 12289 32064 12353 32068
rect 16488 32124 16552 32128
rect 16488 32068 16492 32124
rect 16492 32068 16548 32124
rect 16548 32068 16552 32124
rect 16488 32064 16552 32068
rect 16568 32124 16632 32128
rect 16568 32068 16572 32124
rect 16572 32068 16628 32124
rect 16628 32068 16632 32124
rect 16568 32064 16632 32068
rect 16648 32124 16712 32128
rect 16648 32068 16652 32124
rect 16652 32068 16708 32124
rect 16708 32068 16712 32124
rect 16648 32064 16712 32068
rect 16728 32124 16792 32128
rect 16728 32068 16732 32124
rect 16732 32068 16788 32124
rect 16788 32068 16792 32124
rect 16728 32064 16792 32068
rect 5390 31580 5454 31584
rect 5390 31524 5394 31580
rect 5394 31524 5450 31580
rect 5450 31524 5454 31580
rect 5390 31520 5454 31524
rect 5470 31580 5534 31584
rect 5470 31524 5474 31580
rect 5474 31524 5530 31580
rect 5530 31524 5534 31580
rect 5470 31520 5534 31524
rect 5550 31580 5614 31584
rect 5550 31524 5554 31580
rect 5554 31524 5610 31580
rect 5610 31524 5614 31580
rect 5550 31520 5614 31524
rect 5630 31580 5694 31584
rect 5630 31524 5634 31580
rect 5634 31524 5690 31580
rect 5690 31524 5694 31580
rect 5630 31520 5694 31524
rect 9829 31580 9893 31584
rect 9829 31524 9833 31580
rect 9833 31524 9889 31580
rect 9889 31524 9893 31580
rect 9829 31520 9893 31524
rect 9909 31580 9973 31584
rect 9909 31524 9913 31580
rect 9913 31524 9969 31580
rect 9969 31524 9973 31580
rect 9909 31520 9973 31524
rect 9989 31580 10053 31584
rect 9989 31524 9993 31580
rect 9993 31524 10049 31580
rect 10049 31524 10053 31580
rect 9989 31520 10053 31524
rect 10069 31580 10133 31584
rect 10069 31524 10073 31580
rect 10073 31524 10129 31580
rect 10129 31524 10133 31580
rect 10069 31520 10133 31524
rect 14268 31580 14332 31584
rect 14268 31524 14272 31580
rect 14272 31524 14328 31580
rect 14328 31524 14332 31580
rect 14268 31520 14332 31524
rect 14348 31580 14412 31584
rect 14348 31524 14352 31580
rect 14352 31524 14408 31580
rect 14408 31524 14412 31580
rect 14348 31520 14412 31524
rect 14428 31580 14492 31584
rect 14428 31524 14432 31580
rect 14432 31524 14488 31580
rect 14488 31524 14492 31580
rect 14428 31520 14492 31524
rect 14508 31580 14572 31584
rect 14508 31524 14512 31580
rect 14512 31524 14568 31580
rect 14568 31524 14572 31580
rect 14508 31520 14572 31524
rect 18707 31580 18771 31584
rect 18707 31524 18711 31580
rect 18711 31524 18767 31580
rect 18767 31524 18771 31580
rect 18707 31520 18771 31524
rect 18787 31580 18851 31584
rect 18787 31524 18791 31580
rect 18791 31524 18847 31580
rect 18847 31524 18851 31580
rect 18787 31520 18851 31524
rect 18867 31580 18931 31584
rect 18867 31524 18871 31580
rect 18871 31524 18927 31580
rect 18927 31524 18931 31580
rect 18867 31520 18931 31524
rect 18947 31580 19011 31584
rect 18947 31524 18951 31580
rect 18951 31524 19007 31580
rect 19007 31524 19011 31580
rect 18947 31520 19011 31524
rect 3171 31036 3235 31040
rect 3171 30980 3175 31036
rect 3175 30980 3231 31036
rect 3231 30980 3235 31036
rect 3171 30976 3235 30980
rect 3251 31036 3315 31040
rect 3251 30980 3255 31036
rect 3255 30980 3311 31036
rect 3311 30980 3315 31036
rect 3251 30976 3315 30980
rect 3331 31036 3395 31040
rect 3331 30980 3335 31036
rect 3335 30980 3391 31036
rect 3391 30980 3395 31036
rect 3331 30976 3395 30980
rect 3411 31036 3475 31040
rect 3411 30980 3415 31036
rect 3415 30980 3471 31036
rect 3471 30980 3475 31036
rect 3411 30976 3475 30980
rect 7610 31036 7674 31040
rect 7610 30980 7614 31036
rect 7614 30980 7670 31036
rect 7670 30980 7674 31036
rect 7610 30976 7674 30980
rect 7690 31036 7754 31040
rect 7690 30980 7694 31036
rect 7694 30980 7750 31036
rect 7750 30980 7754 31036
rect 7690 30976 7754 30980
rect 7770 31036 7834 31040
rect 7770 30980 7774 31036
rect 7774 30980 7830 31036
rect 7830 30980 7834 31036
rect 7770 30976 7834 30980
rect 7850 31036 7914 31040
rect 7850 30980 7854 31036
rect 7854 30980 7910 31036
rect 7910 30980 7914 31036
rect 7850 30976 7914 30980
rect 12049 31036 12113 31040
rect 12049 30980 12053 31036
rect 12053 30980 12109 31036
rect 12109 30980 12113 31036
rect 12049 30976 12113 30980
rect 12129 31036 12193 31040
rect 12129 30980 12133 31036
rect 12133 30980 12189 31036
rect 12189 30980 12193 31036
rect 12129 30976 12193 30980
rect 12209 31036 12273 31040
rect 12209 30980 12213 31036
rect 12213 30980 12269 31036
rect 12269 30980 12273 31036
rect 12209 30976 12273 30980
rect 12289 31036 12353 31040
rect 12289 30980 12293 31036
rect 12293 30980 12349 31036
rect 12349 30980 12353 31036
rect 12289 30976 12353 30980
rect 16488 31036 16552 31040
rect 16488 30980 16492 31036
rect 16492 30980 16548 31036
rect 16548 30980 16552 31036
rect 16488 30976 16552 30980
rect 16568 31036 16632 31040
rect 16568 30980 16572 31036
rect 16572 30980 16628 31036
rect 16628 30980 16632 31036
rect 16568 30976 16632 30980
rect 16648 31036 16712 31040
rect 16648 30980 16652 31036
rect 16652 30980 16708 31036
rect 16708 30980 16712 31036
rect 16648 30976 16712 30980
rect 16728 31036 16792 31040
rect 16728 30980 16732 31036
rect 16732 30980 16788 31036
rect 16788 30980 16792 31036
rect 16728 30976 16792 30980
rect 5390 30492 5454 30496
rect 5390 30436 5394 30492
rect 5394 30436 5450 30492
rect 5450 30436 5454 30492
rect 5390 30432 5454 30436
rect 5470 30492 5534 30496
rect 5470 30436 5474 30492
rect 5474 30436 5530 30492
rect 5530 30436 5534 30492
rect 5470 30432 5534 30436
rect 5550 30492 5614 30496
rect 5550 30436 5554 30492
rect 5554 30436 5610 30492
rect 5610 30436 5614 30492
rect 5550 30432 5614 30436
rect 5630 30492 5694 30496
rect 5630 30436 5634 30492
rect 5634 30436 5690 30492
rect 5690 30436 5694 30492
rect 5630 30432 5694 30436
rect 9829 30492 9893 30496
rect 9829 30436 9833 30492
rect 9833 30436 9889 30492
rect 9889 30436 9893 30492
rect 9829 30432 9893 30436
rect 9909 30492 9973 30496
rect 9909 30436 9913 30492
rect 9913 30436 9969 30492
rect 9969 30436 9973 30492
rect 9909 30432 9973 30436
rect 9989 30492 10053 30496
rect 9989 30436 9993 30492
rect 9993 30436 10049 30492
rect 10049 30436 10053 30492
rect 9989 30432 10053 30436
rect 10069 30492 10133 30496
rect 10069 30436 10073 30492
rect 10073 30436 10129 30492
rect 10129 30436 10133 30492
rect 10069 30432 10133 30436
rect 14268 30492 14332 30496
rect 14268 30436 14272 30492
rect 14272 30436 14328 30492
rect 14328 30436 14332 30492
rect 14268 30432 14332 30436
rect 14348 30492 14412 30496
rect 14348 30436 14352 30492
rect 14352 30436 14408 30492
rect 14408 30436 14412 30492
rect 14348 30432 14412 30436
rect 14428 30492 14492 30496
rect 14428 30436 14432 30492
rect 14432 30436 14488 30492
rect 14488 30436 14492 30492
rect 14428 30432 14492 30436
rect 14508 30492 14572 30496
rect 14508 30436 14512 30492
rect 14512 30436 14568 30492
rect 14568 30436 14572 30492
rect 14508 30432 14572 30436
rect 18707 30492 18771 30496
rect 18707 30436 18711 30492
rect 18711 30436 18767 30492
rect 18767 30436 18771 30492
rect 18707 30432 18771 30436
rect 18787 30492 18851 30496
rect 18787 30436 18791 30492
rect 18791 30436 18847 30492
rect 18847 30436 18851 30492
rect 18787 30432 18851 30436
rect 18867 30492 18931 30496
rect 18867 30436 18871 30492
rect 18871 30436 18927 30492
rect 18927 30436 18931 30492
rect 18867 30432 18931 30436
rect 18947 30492 19011 30496
rect 18947 30436 18951 30492
rect 18951 30436 19007 30492
rect 19007 30436 19011 30492
rect 18947 30432 19011 30436
rect 4660 30424 4724 30428
rect 4660 30368 4710 30424
rect 4710 30368 4724 30424
rect 4660 30364 4724 30368
rect 3171 29948 3235 29952
rect 3171 29892 3175 29948
rect 3175 29892 3231 29948
rect 3231 29892 3235 29948
rect 3171 29888 3235 29892
rect 3251 29948 3315 29952
rect 3251 29892 3255 29948
rect 3255 29892 3311 29948
rect 3311 29892 3315 29948
rect 3251 29888 3315 29892
rect 3331 29948 3395 29952
rect 3331 29892 3335 29948
rect 3335 29892 3391 29948
rect 3391 29892 3395 29948
rect 3331 29888 3395 29892
rect 3411 29948 3475 29952
rect 3411 29892 3415 29948
rect 3415 29892 3471 29948
rect 3471 29892 3475 29948
rect 3411 29888 3475 29892
rect 7610 29948 7674 29952
rect 7610 29892 7614 29948
rect 7614 29892 7670 29948
rect 7670 29892 7674 29948
rect 7610 29888 7674 29892
rect 7690 29948 7754 29952
rect 7690 29892 7694 29948
rect 7694 29892 7750 29948
rect 7750 29892 7754 29948
rect 7690 29888 7754 29892
rect 7770 29948 7834 29952
rect 7770 29892 7774 29948
rect 7774 29892 7830 29948
rect 7830 29892 7834 29948
rect 7770 29888 7834 29892
rect 7850 29948 7914 29952
rect 7850 29892 7854 29948
rect 7854 29892 7910 29948
rect 7910 29892 7914 29948
rect 7850 29888 7914 29892
rect 12049 29948 12113 29952
rect 12049 29892 12053 29948
rect 12053 29892 12109 29948
rect 12109 29892 12113 29948
rect 12049 29888 12113 29892
rect 12129 29948 12193 29952
rect 12129 29892 12133 29948
rect 12133 29892 12189 29948
rect 12189 29892 12193 29948
rect 12129 29888 12193 29892
rect 12209 29948 12273 29952
rect 12209 29892 12213 29948
rect 12213 29892 12269 29948
rect 12269 29892 12273 29948
rect 12209 29888 12273 29892
rect 12289 29948 12353 29952
rect 12289 29892 12293 29948
rect 12293 29892 12349 29948
rect 12349 29892 12353 29948
rect 12289 29888 12353 29892
rect 16488 29948 16552 29952
rect 16488 29892 16492 29948
rect 16492 29892 16548 29948
rect 16548 29892 16552 29948
rect 16488 29888 16552 29892
rect 16568 29948 16632 29952
rect 16568 29892 16572 29948
rect 16572 29892 16628 29948
rect 16628 29892 16632 29948
rect 16568 29888 16632 29892
rect 16648 29948 16712 29952
rect 16648 29892 16652 29948
rect 16652 29892 16708 29948
rect 16708 29892 16712 29948
rect 16648 29888 16712 29892
rect 16728 29948 16792 29952
rect 16728 29892 16732 29948
rect 16732 29892 16788 29948
rect 16788 29892 16792 29948
rect 16728 29888 16792 29892
rect 5390 29404 5454 29408
rect 5390 29348 5394 29404
rect 5394 29348 5450 29404
rect 5450 29348 5454 29404
rect 5390 29344 5454 29348
rect 5470 29404 5534 29408
rect 5470 29348 5474 29404
rect 5474 29348 5530 29404
rect 5530 29348 5534 29404
rect 5470 29344 5534 29348
rect 5550 29404 5614 29408
rect 5550 29348 5554 29404
rect 5554 29348 5610 29404
rect 5610 29348 5614 29404
rect 5550 29344 5614 29348
rect 5630 29404 5694 29408
rect 5630 29348 5634 29404
rect 5634 29348 5690 29404
rect 5690 29348 5694 29404
rect 5630 29344 5694 29348
rect 9829 29404 9893 29408
rect 9829 29348 9833 29404
rect 9833 29348 9889 29404
rect 9889 29348 9893 29404
rect 9829 29344 9893 29348
rect 9909 29404 9973 29408
rect 9909 29348 9913 29404
rect 9913 29348 9969 29404
rect 9969 29348 9973 29404
rect 9909 29344 9973 29348
rect 9989 29404 10053 29408
rect 9989 29348 9993 29404
rect 9993 29348 10049 29404
rect 10049 29348 10053 29404
rect 9989 29344 10053 29348
rect 10069 29404 10133 29408
rect 10069 29348 10073 29404
rect 10073 29348 10129 29404
rect 10129 29348 10133 29404
rect 10069 29344 10133 29348
rect 14268 29404 14332 29408
rect 14268 29348 14272 29404
rect 14272 29348 14328 29404
rect 14328 29348 14332 29404
rect 14268 29344 14332 29348
rect 14348 29404 14412 29408
rect 14348 29348 14352 29404
rect 14352 29348 14408 29404
rect 14408 29348 14412 29404
rect 14348 29344 14412 29348
rect 14428 29404 14492 29408
rect 14428 29348 14432 29404
rect 14432 29348 14488 29404
rect 14488 29348 14492 29404
rect 14428 29344 14492 29348
rect 14508 29404 14572 29408
rect 14508 29348 14512 29404
rect 14512 29348 14568 29404
rect 14568 29348 14572 29404
rect 14508 29344 14572 29348
rect 18707 29404 18771 29408
rect 18707 29348 18711 29404
rect 18711 29348 18767 29404
rect 18767 29348 18771 29404
rect 18707 29344 18771 29348
rect 18787 29404 18851 29408
rect 18787 29348 18791 29404
rect 18791 29348 18847 29404
rect 18847 29348 18851 29404
rect 18787 29344 18851 29348
rect 18867 29404 18931 29408
rect 18867 29348 18871 29404
rect 18871 29348 18927 29404
rect 18927 29348 18931 29404
rect 18867 29344 18931 29348
rect 18947 29404 19011 29408
rect 18947 29348 18951 29404
rect 18951 29348 19007 29404
rect 19007 29348 19011 29404
rect 18947 29344 19011 29348
rect 8156 29064 8220 29068
rect 8156 29008 8170 29064
rect 8170 29008 8220 29064
rect 8156 29004 8220 29008
rect 3171 28860 3235 28864
rect 3171 28804 3175 28860
rect 3175 28804 3231 28860
rect 3231 28804 3235 28860
rect 3171 28800 3235 28804
rect 3251 28860 3315 28864
rect 3251 28804 3255 28860
rect 3255 28804 3311 28860
rect 3311 28804 3315 28860
rect 3251 28800 3315 28804
rect 3331 28860 3395 28864
rect 3331 28804 3335 28860
rect 3335 28804 3391 28860
rect 3391 28804 3395 28860
rect 3331 28800 3395 28804
rect 3411 28860 3475 28864
rect 3411 28804 3415 28860
rect 3415 28804 3471 28860
rect 3471 28804 3475 28860
rect 3411 28800 3475 28804
rect 7610 28860 7674 28864
rect 7610 28804 7614 28860
rect 7614 28804 7670 28860
rect 7670 28804 7674 28860
rect 7610 28800 7674 28804
rect 7690 28860 7754 28864
rect 7690 28804 7694 28860
rect 7694 28804 7750 28860
rect 7750 28804 7754 28860
rect 7690 28800 7754 28804
rect 7770 28860 7834 28864
rect 7770 28804 7774 28860
rect 7774 28804 7830 28860
rect 7830 28804 7834 28860
rect 7770 28800 7834 28804
rect 7850 28860 7914 28864
rect 7850 28804 7854 28860
rect 7854 28804 7910 28860
rect 7910 28804 7914 28860
rect 7850 28800 7914 28804
rect 12049 28860 12113 28864
rect 12049 28804 12053 28860
rect 12053 28804 12109 28860
rect 12109 28804 12113 28860
rect 12049 28800 12113 28804
rect 12129 28860 12193 28864
rect 12129 28804 12133 28860
rect 12133 28804 12189 28860
rect 12189 28804 12193 28860
rect 12129 28800 12193 28804
rect 12209 28860 12273 28864
rect 12209 28804 12213 28860
rect 12213 28804 12269 28860
rect 12269 28804 12273 28860
rect 12209 28800 12273 28804
rect 12289 28860 12353 28864
rect 12289 28804 12293 28860
rect 12293 28804 12349 28860
rect 12349 28804 12353 28860
rect 12289 28800 12353 28804
rect 16488 28860 16552 28864
rect 16488 28804 16492 28860
rect 16492 28804 16548 28860
rect 16548 28804 16552 28860
rect 16488 28800 16552 28804
rect 16568 28860 16632 28864
rect 16568 28804 16572 28860
rect 16572 28804 16628 28860
rect 16628 28804 16632 28860
rect 16568 28800 16632 28804
rect 16648 28860 16712 28864
rect 16648 28804 16652 28860
rect 16652 28804 16708 28860
rect 16708 28804 16712 28860
rect 16648 28800 16712 28804
rect 16728 28860 16792 28864
rect 16728 28804 16732 28860
rect 16732 28804 16788 28860
rect 16788 28804 16792 28860
rect 16728 28800 16792 28804
rect 5390 28316 5454 28320
rect 5390 28260 5394 28316
rect 5394 28260 5450 28316
rect 5450 28260 5454 28316
rect 5390 28256 5454 28260
rect 5470 28316 5534 28320
rect 5470 28260 5474 28316
rect 5474 28260 5530 28316
rect 5530 28260 5534 28316
rect 5470 28256 5534 28260
rect 5550 28316 5614 28320
rect 5550 28260 5554 28316
rect 5554 28260 5610 28316
rect 5610 28260 5614 28316
rect 5550 28256 5614 28260
rect 5630 28316 5694 28320
rect 5630 28260 5634 28316
rect 5634 28260 5690 28316
rect 5690 28260 5694 28316
rect 5630 28256 5694 28260
rect 9829 28316 9893 28320
rect 9829 28260 9833 28316
rect 9833 28260 9889 28316
rect 9889 28260 9893 28316
rect 9829 28256 9893 28260
rect 9909 28316 9973 28320
rect 9909 28260 9913 28316
rect 9913 28260 9969 28316
rect 9969 28260 9973 28316
rect 9909 28256 9973 28260
rect 9989 28316 10053 28320
rect 9989 28260 9993 28316
rect 9993 28260 10049 28316
rect 10049 28260 10053 28316
rect 9989 28256 10053 28260
rect 10069 28316 10133 28320
rect 10069 28260 10073 28316
rect 10073 28260 10129 28316
rect 10129 28260 10133 28316
rect 10069 28256 10133 28260
rect 14268 28316 14332 28320
rect 14268 28260 14272 28316
rect 14272 28260 14328 28316
rect 14328 28260 14332 28316
rect 14268 28256 14332 28260
rect 14348 28316 14412 28320
rect 14348 28260 14352 28316
rect 14352 28260 14408 28316
rect 14408 28260 14412 28316
rect 14348 28256 14412 28260
rect 14428 28316 14492 28320
rect 14428 28260 14432 28316
rect 14432 28260 14488 28316
rect 14488 28260 14492 28316
rect 14428 28256 14492 28260
rect 14508 28316 14572 28320
rect 14508 28260 14512 28316
rect 14512 28260 14568 28316
rect 14568 28260 14572 28316
rect 14508 28256 14572 28260
rect 18707 28316 18771 28320
rect 18707 28260 18711 28316
rect 18711 28260 18767 28316
rect 18767 28260 18771 28316
rect 18707 28256 18771 28260
rect 18787 28316 18851 28320
rect 18787 28260 18791 28316
rect 18791 28260 18847 28316
rect 18847 28260 18851 28316
rect 18787 28256 18851 28260
rect 18867 28316 18931 28320
rect 18867 28260 18871 28316
rect 18871 28260 18927 28316
rect 18927 28260 18931 28316
rect 18867 28256 18931 28260
rect 18947 28316 19011 28320
rect 18947 28260 18951 28316
rect 18951 28260 19007 28316
rect 19007 28260 19011 28316
rect 18947 28256 19011 28260
rect 3171 27772 3235 27776
rect 3171 27716 3175 27772
rect 3175 27716 3231 27772
rect 3231 27716 3235 27772
rect 3171 27712 3235 27716
rect 3251 27772 3315 27776
rect 3251 27716 3255 27772
rect 3255 27716 3311 27772
rect 3311 27716 3315 27772
rect 3251 27712 3315 27716
rect 3331 27772 3395 27776
rect 3331 27716 3335 27772
rect 3335 27716 3391 27772
rect 3391 27716 3395 27772
rect 3331 27712 3395 27716
rect 3411 27772 3475 27776
rect 3411 27716 3415 27772
rect 3415 27716 3471 27772
rect 3471 27716 3475 27772
rect 3411 27712 3475 27716
rect 7610 27772 7674 27776
rect 7610 27716 7614 27772
rect 7614 27716 7670 27772
rect 7670 27716 7674 27772
rect 7610 27712 7674 27716
rect 7690 27772 7754 27776
rect 7690 27716 7694 27772
rect 7694 27716 7750 27772
rect 7750 27716 7754 27772
rect 7690 27712 7754 27716
rect 7770 27772 7834 27776
rect 7770 27716 7774 27772
rect 7774 27716 7830 27772
rect 7830 27716 7834 27772
rect 7770 27712 7834 27716
rect 7850 27772 7914 27776
rect 7850 27716 7854 27772
rect 7854 27716 7910 27772
rect 7910 27716 7914 27772
rect 7850 27712 7914 27716
rect 12049 27772 12113 27776
rect 12049 27716 12053 27772
rect 12053 27716 12109 27772
rect 12109 27716 12113 27772
rect 12049 27712 12113 27716
rect 12129 27772 12193 27776
rect 12129 27716 12133 27772
rect 12133 27716 12189 27772
rect 12189 27716 12193 27772
rect 12129 27712 12193 27716
rect 12209 27772 12273 27776
rect 12209 27716 12213 27772
rect 12213 27716 12269 27772
rect 12269 27716 12273 27772
rect 12209 27712 12273 27716
rect 12289 27772 12353 27776
rect 12289 27716 12293 27772
rect 12293 27716 12349 27772
rect 12349 27716 12353 27772
rect 12289 27712 12353 27716
rect 16488 27772 16552 27776
rect 16488 27716 16492 27772
rect 16492 27716 16548 27772
rect 16548 27716 16552 27772
rect 16488 27712 16552 27716
rect 16568 27772 16632 27776
rect 16568 27716 16572 27772
rect 16572 27716 16628 27772
rect 16628 27716 16632 27772
rect 16568 27712 16632 27716
rect 16648 27772 16712 27776
rect 16648 27716 16652 27772
rect 16652 27716 16708 27772
rect 16708 27716 16712 27772
rect 16648 27712 16712 27716
rect 16728 27772 16792 27776
rect 16728 27716 16732 27772
rect 16732 27716 16788 27772
rect 16788 27716 16792 27772
rect 16728 27712 16792 27716
rect 4292 27704 4356 27708
rect 4292 27648 4306 27704
rect 4306 27648 4356 27704
rect 4292 27644 4356 27648
rect 5390 27228 5454 27232
rect 5390 27172 5394 27228
rect 5394 27172 5450 27228
rect 5450 27172 5454 27228
rect 5390 27168 5454 27172
rect 5470 27228 5534 27232
rect 5470 27172 5474 27228
rect 5474 27172 5530 27228
rect 5530 27172 5534 27228
rect 5470 27168 5534 27172
rect 5550 27228 5614 27232
rect 5550 27172 5554 27228
rect 5554 27172 5610 27228
rect 5610 27172 5614 27228
rect 5550 27168 5614 27172
rect 5630 27228 5694 27232
rect 5630 27172 5634 27228
rect 5634 27172 5690 27228
rect 5690 27172 5694 27228
rect 5630 27168 5694 27172
rect 9829 27228 9893 27232
rect 9829 27172 9833 27228
rect 9833 27172 9889 27228
rect 9889 27172 9893 27228
rect 9829 27168 9893 27172
rect 9909 27228 9973 27232
rect 9909 27172 9913 27228
rect 9913 27172 9969 27228
rect 9969 27172 9973 27228
rect 9909 27168 9973 27172
rect 9989 27228 10053 27232
rect 9989 27172 9993 27228
rect 9993 27172 10049 27228
rect 10049 27172 10053 27228
rect 9989 27168 10053 27172
rect 10069 27228 10133 27232
rect 10069 27172 10073 27228
rect 10073 27172 10129 27228
rect 10129 27172 10133 27228
rect 10069 27168 10133 27172
rect 14268 27228 14332 27232
rect 14268 27172 14272 27228
rect 14272 27172 14328 27228
rect 14328 27172 14332 27228
rect 14268 27168 14332 27172
rect 14348 27228 14412 27232
rect 14348 27172 14352 27228
rect 14352 27172 14408 27228
rect 14408 27172 14412 27228
rect 14348 27168 14412 27172
rect 14428 27228 14492 27232
rect 14428 27172 14432 27228
rect 14432 27172 14488 27228
rect 14488 27172 14492 27228
rect 14428 27168 14492 27172
rect 14508 27228 14572 27232
rect 14508 27172 14512 27228
rect 14512 27172 14568 27228
rect 14568 27172 14572 27228
rect 14508 27168 14572 27172
rect 18707 27228 18771 27232
rect 18707 27172 18711 27228
rect 18711 27172 18767 27228
rect 18767 27172 18771 27228
rect 18707 27168 18771 27172
rect 18787 27228 18851 27232
rect 18787 27172 18791 27228
rect 18791 27172 18847 27228
rect 18847 27172 18851 27228
rect 18787 27168 18851 27172
rect 18867 27228 18931 27232
rect 18867 27172 18871 27228
rect 18871 27172 18927 27228
rect 18927 27172 18931 27228
rect 18867 27168 18931 27172
rect 18947 27228 19011 27232
rect 18947 27172 18951 27228
rect 18951 27172 19007 27228
rect 19007 27172 19011 27228
rect 18947 27168 19011 27172
rect 7420 27160 7484 27164
rect 7420 27104 7470 27160
rect 7470 27104 7484 27160
rect 7420 27100 7484 27104
rect 3171 26684 3235 26688
rect 3171 26628 3175 26684
rect 3175 26628 3231 26684
rect 3231 26628 3235 26684
rect 3171 26624 3235 26628
rect 3251 26684 3315 26688
rect 3251 26628 3255 26684
rect 3255 26628 3311 26684
rect 3311 26628 3315 26684
rect 3251 26624 3315 26628
rect 3331 26684 3395 26688
rect 3331 26628 3335 26684
rect 3335 26628 3391 26684
rect 3391 26628 3395 26684
rect 3331 26624 3395 26628
rect 3411 26684 3475 26688
rect 3411 26628 3415 26684
rect 3415 26628 3471 26684
rect 3471 26628 3475 26684
rect 3411 26624 3475 26628
rect 7610 26684 7674 26688
rect 7610 26628 7614 26684
rect 7614 26628 7670 26684
rect 7670 26628 7674 26684
rect 7610 26624 7674 26628
rect 7690 26684 7754 26688
rect 7690 26628 7694 26684
rect 7694 26628 7750 26684
rect 7750 26628 7754 26684
rect 7690 26624 7754 26628
rect 7770 26684 7834 26688
rect 7770 26628 7774 26684
rect 7774 26628 7830 26684
rect 7830 26628 7834 26684
rect 7770 26624 7834 26628
rect 7850 26684 7914 26688
rect 7850 26628 7854 26684
rect 7854 26628 7910 26684
rect 7910 26628 7914 26684
rect 7850 26624 7914 26628
rect 12049 26684 12113 26688
rect 12049 26628 12053 26684
rect 12053 26628 12109 26684
rect 12109 26628 12113 26684
rect 12049 26624 12113 26628
rect 12129 26684 12193 26688
rect 12129 26628 12133 26684
rect 12133 26628 12189 26684
rect 12189 26628 12193 26684
rect 12129 26624 12193 26628
rect 12209 26684 12273 26688
rect 12209 26628 12213 26684
rect 12213 26628 12269 26684
rect 12269 26628 12273 26684
rect 12209 26624 12273 26628
rect 12289 26684 12353 26688
rect 12289 26628 12293 26684
rect 12293 26628 12349 26684
rect 12349 26628 12353 26684
rect 12289 26624 12353 26628
rect 16488 26684 16552 26688
rect 16488 26628 16492 26684
rect 16492 26628 16548 26684
rect 16548 26628 16552 26684
rect 16488 26624 16552 26628
rect 16568 26684 16632 26688
rect 16568 26628 16572 26684
rect 16572 26628 16628 26684
rect 16628 26628 16632 26684
rect 16568 26624 16632 26628
rect 16648 26684 16712 26688
rect 16648 26628 16652 26684
rect 16652 26628 16708 26684
rect 16708 26628 16712 26684
rect 16648 26624 16712 26628
rect 16728 26684 16792 26688
rect 16728 26628 16732 26684
rect 16732 26628 16788 26684
rect 16788 26628 16792 26684
rect 16728 26624 16792 26628
rect 1900 26556 1964 26620
rect 6684 26284 6748 26348
rect 5390 26140 5454 26144
rect 5390 26084 5394 26140
rect 5394 26084 5450 26140
rect 5450 26084 5454 26140
rect 5390 26080 5454 26084
rect 5470 26140 5534 26144
rect 5470 26084 5474 26140
rect 5474 26084 5530 26140
rect 5530 26084 5534 26140
rect 5470 26080 5534 26084
rect 5550 26140 5614 26144
rect 5550 26084 5554 26140
rect 5554 26084 5610 26140
rect 5610 26084 5614 26140
rect 5550 26080 5614 26084
rect 5630 26140 5694 26144
rect 5630 26084 5634 26140
rect 5634 26084 5690 26140
rect 5690 26084 5694 26140
rect 5630 26080 5694 26084
rect 9829 26140 9893 26144
rect 9829 26084 9833 26140
rect 9833 26084 9889 26140
rect 9889 26084 9893 26140
rect 9829 26080 9893 26084
rect 9909 26140 9973 26144
rect 9909 26084 9913 26140
rect 9913 26084 9969 26140
rect 9969 26084 9973 26140
rect 9909 26080 9973 26084
rect 9989 26140 10053 26144
rect 9989 26084 9993 26140
rect 9993 26084 10049 26140
rect 10049 26084 10053 26140
rect 9989 26080 10053 26084
rect 10069 26140 10133 26144
rect 10069 26084 10073 26140
rect 10073 26084 10129 26140
rect 10129 26084 10133 26140
rect 10069 26080 10133 26084
rect 14268 26140 14332 26144
rect 14268 26084 14272 26140
rect 14272 26084 14328 26140
rect 14328 26084 14332 26140
rect 14268 26080 14332 26084
rect 14348 26140 14412 26144
rect 14348 26084 14352 26140
rect 14352 26084 14408 26140
rect 14408 26084 14412 26140
rect 14348 26080 14412 26084
rect 14428 26140 14492 26144
rect 14428 26084 14432 26140
rect 14432 26084 14488 26140
rect 14488 26084 14492 26140
rect 14428 26080 14492 26084
rect 14508 26140 14572 26144
rect 14508 26084 14512 26140
rect 14512 26084 14568 26140
rect 14568 26084 14572 26140
rect 14508 26080 14572 26084
rect 18707 26140 18771 26144
rect 18707 26084 18711 26140
rect 18711 26084 18767 26140
rect 18767 26084 18771 26140
rect 18707 26080 18771 26084
rect 18787 26140 18851 26144
rect 18787 26084 18791 26140
rect 18791 26084 18847 26140
rect 18847 26084 18851 26140
rect 18787 26080 18851 26084
rect 18867 26140 18931 26144
rect 18867 26084 18871 26140
rect 18871 26084 18927 26140
rect 18927 26084 18931 26140
rect 18867 26080 18931 26084
rect 18947 26140 19011 26144
rect 18947 26084 18951 26140
rect 18951 26084 19007 26140
rect 19007 26084 19011 26140
rect 18947 26080 19011 26084
rect 3171 25596 3235 25600
rect 3171 25540 3175 25596
rect 3175 25540 3231 25596
rect 3231 25540 3235 25596
rect 3171 25536 3235 25540
rect 3251 25596 3315 25600
rect 3251 25540 3255 25596
rect 3255 25540 3311 25596
rect 3311 25540 3315 25596
rect 3251 25536 3315 25540
rect 3331 25596 3395 25600
rect 3331 25540 3335 25596
rect 3335 25540 3391 25596
rect 3391 25540 3395 25596
rect 3331 25536 3395 25540
rect 3411 25596 3475 25600
rect 3411 25540 3415 25596
rect 3415 25540 3471 25596
rect 3471 25540 3475 25596
rect 3411 25536 3475 25540
rect 7610 25596 7674 25600
rect 7610 25540 7614 25596
rect 7614 25540 7670 25596
rect 7670 25540 7674 25596
rect 7610 25536 7674 25540
rect 7690 25596 7754 25600
rect 7690 25540 7694 25596
rect 7694 25540 7750 25596
rect 7750 25540 7754 25596
rect 7690 25536 7754 25540
rect 7770 25596 7834 25600
rect 7770 25540 7774 25596
rect 7774 25540 7830 25596
rect 7830 25540 7834 25596
rect 7770 25536 7834 25540
rect 7850 25596 7914 25600
rect 7850 25540 7854 25596
rect 7854 25540 7910 25596
rect 7910 25540 7914 25596
rect 7850 25536 7914 25540
rect 12049 25596 12113 25600
rect 12049 25540 12053 25596
rect 12053 25540 12109 25596
rect 12109 25540 12113 25596
rect 12049 25536 12113 25540
rect 12129 25596 12193 25600
rect 12129 25540 12133 25596
rect 12133 25540 12189 25596
rect 12189 25540 12193 25596
rect 12129 25536 12193 25540
rect 12209 25596 12273 25600
rect 12209 25540 12213 25596
rect 12213 25540 12269 25596
rect 12269 25540 12273 25596
rect 12209 25536 12273 25540
rect 12289 25596 12353 25600
rect 12289 25540 12293 25596
rect 12293 25540 12349 25596
rect 12349 25540 12353 25596
rect 12289 25536 12353 25540
rect 16488 25596 16552 25600
rect 16488 25540 16492 25596
rect 16492 25540 16548 25596
rect 16548 25540 16552 25596
rect 16488 25536 16552 25540
rect 16568 25596 16632 25600
rect 16568 25540 16572 25596
rect 16572 25540 16628 25596
rect 16628 25540 16632 25596
rect 16568 25536 16632 25540
rect 16648 25596 16712 25600
rect 16648 25540 16652 25596
rect 16652 25540 16708 25596
rect 16708 25540 16712 25596
rect 16648 25536 16712 25540
rect 16728 25596 16792 25600
rect 16728 25540 16732 25596
rect 16732 25540 16788 25596
rect 16788 25540 16792 25596
rect 16728 25536 16792 25540
rect 4844 25196 4908 25260
rect 5390 25052 5454 25056
rect 5390 24996 5394 25052
rect 5394 24996 5450 25052
rect 5450 24996 5454 25052
rect 5390 24992 5454 24996
rect 5470 25052 5534 25056
rect 5470 24996 5474 25052
rect 5474 24996 5530 25052
rect 5530 24996 5534 25052
rect 5470 24992 5534 24996
rect 5550 25052 5614 25056
rect 5550 24996 5554 25052
rect 5554 24996 5610 25052
rect 5610 24996 5614 25052
rect 5550 24992 5614 24996
rect 5630 25052 5694 25056
rect 5630 24996 5634 25052
rect 5634 24996 5690 25052
rect 5690 24996 5694 25052
rect 5630 24992 5694 24996
rect 9829 25052 9893 25056
rect 9829 24996 9833 25052
rect 9833 24996 9889 25052
rect 9889 24996 9893 25052
rect 9829 24992 9893 24996
rect 9909 25052 9973 25056
rect 9909 24996 9913 25052
rect 9913 24996 9969 25052
rect 9969 24996 9973 25052
rect 9909 24992 9973 24996
rect 9989 25052 10053 25056
rect 9989 24996 9993 25052
rect 9993 24996 10049 25052
rect 10049 24996 10053 25052
rect 9989 24992 10053 24996
rect 10069 25052 10133 25056
rect 10069 24996 10073 25052
rect 10073 24996 10129 25052
rect 10129 24996 10133 25052
rect 10069 24992 10133 24996
rect 14268 25052 14332 25056
rect 14268 24996 14272 25052
rect 14272 24996 14328 25052
rect 14328 24996 14332 25052
rect 14268 24992 14332 24996
rect 14348 25052 14412 25056
rect 14348 24996 14352 25052
rect 14352 24996 14408 25052
rect 14408 24996 14412 25052
rect 14348 24992 14412 24996
rect 14428 25052 14492 25056
rect 14428 24996 14432 25052
rect 14432 24996 14488 25052
rect 14488 24996 14492 25052
rect 14428 24992 14492 24996
rect 14508 25052 14572 25056
rect 14508 24996 14512 25052
rect 14512 24996 14568 25052
rect 14568 24996 14572 25052
rect 14508 24992 14572 24996
rect 18707 25052 18771 25056
rect 18707 24996 18711 25052
rect 18711 24996 18767 25052
rect 18767 24996 18771 25052
rect 18707 24992 18771 24996
rect 18787 25052 18851 25056
rect 18787 24996 18791 25052
rect 18791 24996 18847 25052
rect 18847 24996 18851 25052
rect 18787 24992 18851 24996
rect 18867 25052 18931 25056
rect 18867 24996 18871 25052
rect 18871 24996 18927 25052
rect 18927 24996 18931 25052
rect 18867 24992 18931 24996
rect 18947 25052 19011 25056
rect 18947 24996 18951 25052
rect 18951 24996 19007 25052
rect 19007 24996 19011 25052
rect 18947 24992 19011 24996
rect 3171 24508 3235 24512
rect 3171 24452 3175 24508
rect 3175 24452 3231 24508
rect 3231 24452 3235 24508
rect 3171 24448 3235 24452
rect 3251 24508 3315 24512
rect 3251 24452 3255 24508
rect 3255 24452 3311 24508
rect 3311 24452 3315 24508
rect 3251 24448 3315 24452
rect 3331 24508 3395 24512
rect 3331 24452 3335 24508
rect 3335 24452 3391 24508
rect 3391 24452 3395 24508
rect 3331 24448 3395 24452
rect 3411 24508 3475 24512
rect 3411 24452 3415 24508
rect 3415 24452 3471 24508
rect 3471 24452 3475 24508
rect 3411 24448 3475 24452
rect 7610 24508 7674 24512
rect 7610 24452 7614 24508
rect 7614 24452 7670 24508
rect 7670 24452 7674 24508
rect 7610 24448 7674 24452
rect 7690 24508 7754 24512
rect 7690 24452 7694 24508
rect 7694 24452 7750 24508
rect 7750 24452 7754 24508
rect 7690 24448 7754 24452
rect 7770 24508 7834 24512
rect 7770 24452 7774 24508
rect 7774 24452 7830 24508
rect 7830 24452 7834 24508
rect 7770 24448 7834 24452
rect 7850 24508 7914 24512
rect 7850 24452 7854 24508
rect 7854 24452 7910 24508
rect 7910 24452 7914 24508
rect 7850 24448 7914 24452
rect 12049 24508 12113 24512
rect 12049 24452 12053 24508
rect 12053 24452 12109 24508
rect 12109 24452 12113 24508
rect 12049 24448 12113 24452
rect 12129 24508 12193 24512
rect 12129 24452 12133 24508
rect 12133 24452 12189 24508
rect 12189 24452 12193 24508
rect 12129 24448 12193 24452
rect 12209 24508 12273 24512
rect 12209 24452 12213 24508
rect 12213 24452 12269 24508
rect 12269 24452 12273 24508
rect 12209 24448 12273 24452
rect 12289 24508 12353 24512
rect 12289 24452 12293 24508
rect 12293 24452 12349 24508
rect 12349 24452 12353 24508
rect 12289 24448 12353 24452
rect 16488 24508 16552 24512
rect 16488 24452 16492 24508
rect 16492 24452 16548 24508
rect 16548 24452 16552 24508
rect 16488 24448 16552 24452
rect 16568 24508 16632 24512
rect 16568 24452 16572 24508
rect 16572 24452 16628 24508
rect 16628 24452 16632 24508
rect 16568 24448 16632 24452
rect 16648 24508 16712 24512
rect 16648 24452 16652 24508
rect 16652 24452 16708 24508
rect 16708 24452 16712 24508
rect 16648 24448 16712 24452
rect 16728 24508 16792 24512
rect 16728 24452 16732 24508
rect 16732 24452 16788 24508
rect 16788 24452 16792 24508
rect 16728 24448 16792 24452
rect 7420 24108 7484 24172
rect 5390 23964 5454 23968
rect 5390 23908 5394 23964
rect 5394 23908 5450 23964
rect 5450 23908 5454 23964
rect 5390 23904 5454 23908
rect 5470 23964 5534 23968
rect 5470 23908 5474 23964
rect 5474 23908 5530 23964
rect 5530 23908 5534 23964
rect 5470 23904 5534 23908
rect 5550 23964 5614 23968
rect 5550 23908 5554 23964
rect 5554 23908 5610 23964
rect 5610 23908 5614 23964
rect 5550 23904 5614 23908
rect 5630 23964 5694 23968
rect 5630 23908 5634 23964
rect 5634 23908 5690 23964
rect 5690 23908 5694 23964
rect 5630 23904 5694 23908
rect 9829 23964 9893 23968
rect 9829 23908 9833 23964
rect 9833 23908 9889 23964
rect 9889 23908 9893 23964
rect 9829 23904 9893 23908
rect 9909 23964 9973 23968
rect 9909 23908 9913 23964
rect 9913 23908 9969 23964
rect 9969 23908 9973 23964
rect 9909 23904 9973 23908
rect 9989 23964 10053 23968
rect 9989 23908 9993 23964
rect 9993 23908 10049 23964
rect 10049 23908 10053 23964
rect 9989 23904 10053 23908
rect 10069 23964 10133 23968
rect 10069 23908 10073 23964
rect 10073 23908 10129 23964
rect 10129 23908 10133 23964
rect 10069 23904 10133 23908
rect 14268 23964 14332 23968
rect 14268 23908 14272 23964
rect 14272 23908 14328 23964
rect 14328 23908 14332 23964
rect 14268 23904 14332 23908
rect 14348 23964 14412 23968
rect 14348 23908 14352 23964
rect 14352 23908 14408 23964
rect 14408 23908 14412 23964
rect 14348 23904 14412 23908
rect 14428 23964 14492 23968
rect 14428 23908 14432 23964
rect 14432 23908 14488 23964
rect 14488 23908 14492 23964
rect 14428 23904 14492 23908
rect 14508 23964 14572 23968
rect 14508 23908 14512 23964
rect 14512 23908 14568 23964
rect 14568 23908 14572 23964
rect 14508 23904 14572 23908
rect 18707 23964 18771 23968
rect 18707 23908 18711 23964
rect 18711 23908 18767 23964
rect 18767 23908 18771 23964
rect 18707 23904 18771 23908
rect 18787 23964 18851 23968
rect 18787 23908 18791 23964
rect 18791 23908 18847 23964
rect 18847 23908 18851 23964
rect 18787 23904 18851 23908
rect 18867 23964 18931 23968
rect 18867 23908 18871 23964
rect 18871 23908 18927 23964
rect 18927 23908 18931 23964
rect 18867 23904 18931 23908
rect 18947 23964 19011 23968
rect 18947 23908 18951 23964
rect 18951 23908 19007 23964
rect 19007 23908 19011 23964
rect 18947 23904 19011 23908
rect 3924 23428 3988 23492
rect 3171 23420 3235 23424
rect 3171 23364 3175 23420
rect 3175 23364 3231 23420
rect 3231 23364 3235 23420
rect 3171 23360 3235 23364
rect 3251 23420 3315 23424
rect 3251 23364 3255 23420
rect 3255 23364 3311 23420
rect 3311 23364 3315 23420
rect 3251 23360 3315 23364
rect 3331 23420 3395 23424
rect 3331 23364 3335 23420
rect 3335 23364 3391 23420
rect 3391 23364 3395 23420
rect 3331 23360 3395 23364
rect 3411 23420 3475 23424
rect 3411 23364 3415 23420
rect 3415 23364 3471 23420
rect 3471 23364 3475 23420
rect 3411 23360 3475 23364
rect 7610 23420 7674 23424
rect 7610 23364 7614 23420
rect 7614 23364 7670 23420
rect 7670 23364 7674 23420
rect 7610 23360 7674 23364
rect 7690 23420 7754 23424
rect 7690 23364 7694 23420
rect 7694 23364 7750 23420
rect 7750 23364 7754 23420
rect 7690 23360 7754 23364
rect 7770 23420 7834 23424
rect 7770 23364 7774 23420
rect 7774 23364 7830 23420
rect 7830 23364 7834 23420
rect 7770 23360 7834 23364
rect 7850 23420 7914 23424
rect 7850 23364 7854 23420
rect 7854 23364 7910 23420
rect 7910 23364 7914 23420
rect 7850 23360 7914 23364
rect 12049 23420 12113 23424
rect 12049 23364 12053 23420
rect 12053 23364 12109 23420
rect 12109 23364 12113 23420
rect 12049 23360 12113 23364
rect 12129 23420 12193 23424
rect 12129 23364 12133 23420
rect 12133 23364 12189 23420
rect 12189 23364 12193 23420
rect 12129 23360 12193 23364
rect 12209 23420 12273 23424
rect 12209 23364 12213 23420
rect 12213 23364 12269 23420
rect 12269 23364 12273 23420
rect 12209 23360 12273 23364
rect 12289 23420 12353 23424
rect 12289 23364 12293 23420
rect 12293 23364 12349 23420
rect 12349 23364 12353 23420
rect 12289 23360 12353 23364
rect 16488 23420 16552 23424
rect 16488 23364 16492 23420
rect 16492 23364 16548 23420
rect 16548 23364 16552 23420
rect 16488 23360 16552 23364
rect 16568 23420 16632 23424
rect 16568 23364 16572 23420
rect 16572 23364 16628 23420
rect 16628 23364 16632 23420
rect 16568 23360 16632 23364
rect 16648 23420 16712 23424
rect 16648 23364 16652 23420
rect 16652 23364 16708 23420
rect 16708 23364 16712 23420
rect 16648 23360 16712 23364
rect 16728 23420 16792 23424
rect 16728 23364 16732 23420
rect 16732 23364 16788 23420
rect 16788 23364 16792 23420
rect 16728 23360 16792 23364
rect 5390 22876 5454 22880
rect 5390 22820 5394 22876
rect 5394 22820 5450 22876
rect 5450 22820 5454 22876
rect 5390 22816 5454 22820
rect 5470 22876 5534 22880
rect 5470 22820 5474 22876
rect 5474 22820 5530 22876
rect 5530 22820 5534 22876
rect 5470 22816 5534 22820
rect 5550 22876 5614 22880
rect 5550 22820 5554 22876
rect 5554 22820 5610 22876
rect 5610 22820 5614 22876
rect 5550 22816 5614 22820
rect 5630 22876 5694 22880
rect 5630 22820 5634 22876
rect 5634 22820 5690 22876
rect 5690 22820 5694 22876
rect 5630 22816 5694 22820
rect 9829 22876 9893 22880
rect 9829 22820 9833 22876
rect 9833 22820 9889 22876
rect 9889 22820 9893 22876
rect 9829 22816 9893 22820
rect 9909 22876 9973 22880
rect 9909 22820 9913 22876
rect 9913 22820 9969 22876
rect 9969 22820 9973 22876
rect 9909 22816 9973 22820
rect 9989 22876 10053 22880
rect 9989 22820 9993 22876
rect 9993 22820 10049 22876
rect 10049 22820 10053 22876
rect 9989 22816 10053 22820
rect 10069 22876 10133 22880
rect 10069 22820 10073 22876
rect 10073 22820 10129 22876
rect 10129 22820 10133 22876
rect 10069 22816 10133 22820
rect 14268 22876 14332 22880
rect 14268 22820 14272 22876
rect 14272 22820 14328 22876
rect 14328 22820 14332 22876
rect 14268 22816 14332 22820
rect 14348 22876 14412 22880
rect 14348 22820 14352 22876
rect 14352 22820 14408 22876
rect 14408 22820 14412 22876
rect 14348 22816 14412 22820
rect 14428 22876 14492 22880
rect 14428 22820 14432 22876
rect 14432 22820 14488 22876
rect 14488 22820 14492 22876
rect 14428 22816 14492 22820
rect 14508 22876 14572 22880
rect 14508 22820 14512 22876
rect 14512 22820 14568 22876
rect 14568 22820 14572 22876
rect 14508 22816 14572 22820
rect 18707 22876 18771 22880
rect 18707 22820 18711 22876
rect 18711 22820 18767 22876
rect 18767 22820 18771 22876
rect 18707 22816 18771 22820
rect 18787 22876 18851 22880
rect 18787 22820 18791 22876
rect 18791 22820 18847 22876
rect 18847 22820 18851 22876
rect 18787 22816 18851 22820
rect 18867 22876 18931 22880
rect 18867 22820 18871 22876
rect 18871 22820 18927 22876
rect 18927 22820 18931 22876
rect 18867 22816 18931 22820
rect 18947 22876 19011 22880
rect 18947 22820 18951 22876
rect 18951 22820 19007 22876
rect 19007 22820 19011 22876
rect 18947 22816 19011 22820
rect 3171 22332 3235 22336
rect 3171 22276 3175 22332
rect 3175 22276 3231 22332
rect 3231 22276 3235 22332
rect 3171 22272 3235 22276
rect 3251 22332 3315 22336
rect 3251 22276 3255 22332
rect 3255 22276 3311 22332
rect 3311 22276 3315 22332
rect 3251 22272 3315 22276
rect 3331 22332 3395 22336
rect 3331 22276 3335 22332
rect 3335 22276 3391 22332
rect 3391 22276 3395 22332
rect 3331 22272 3395 22276
rect 3411 22332 3475 22336
rect 3411 22276 3415 22332
rect 3415 22276 3471 22332
rect 3471 22276 3475 22332
rect 3411 22272 3475 22276
rect 7610 22332 7674 22336
rect 7610 22276 7614 22332
rect 7614 22276 7670 22332
rect 7670 22276 7674 22332
rect 7610 22272 7674 22276
rect 7690 22332 7754 22336
rect 7690 22276 7694 22332
rect 7694 22276 7750 22332
rect 7750 22276 7754 22332
rect 7690 22272 7754 22276
rect 7770 22332 7834 22336
rect 7770 22276 7774 22332
rect 7774 22276 7830 22332
rect 7830 22276 7834 22332
rect 7770 22272 7834 22276
rect 7850 22332 7914 22336
rect 7850 22276 7854 22332
rect 7854 22276 7910 22332
rect 7910 22276 7914 22332
rect 7850 22272 7914 22276
rect 12049 22332 12113 22336
rect 12049 22276 12053 22332
rect 12053 22276 12109 22332
rect 12109 22276 12113 22332
rect 12049 22272 12113 22276
rect 12129 22332 12193 22336
rect 12129 22276 12133 22332
rect 12133 22276 12189 22332
rect 12189 22276 12193 22332
rect 12129 22272 12193 22276
rect 12209 22332 12273 22336
rect 12209 22276 12213 22332
rect 12213 22276 12269 22332
rect 12269 22276 12273 22332
rect 12209 22272 12273 22276
rect 12289 22332 12353 22336
rect 12289 22276 12293 22332
rect 12293 22276 12349 22332
rect 12349 22276 12353 22332
rect 12289 22272 12353 22276
rect 16488 22332 16552 22336
rect 16488 22276 16492 22332
rect 16492 22276 16548 22332
rect 16548 22276 16552 22332
rect 16488 22272 16552 22276
rect 16568 22332 16632 22336
rect 16568 22276 16572 22332
rect 16572 22276 16628 22332
rect 16628 22276 16632 22332
rect 16568 22272 16632 22276
rect 16648 22332 16712 22336
rect 16648 22276 16652 22332
rect 16652 22276 16708 22332
rect 16708 22276 16712 22332
rect 16648 22272 16712 22276
rect 16728 22332 16792 22336
rect 16728 22276 16732 22332
rect 16732 22276 16788 22332
rect 16788 22276 16792 22332
rect 16728 22272 16792 22276
rect 5390 21788 5454 21792
rect 5390 21732 5394 21788
rect 5394 21732 5450 21788
rect 5450 21732 5454 21788
rect 5390 21728 5454 21732
rect 5470 21788 5534 21792
rect 5470 21732 5474 21788
rect 5474 21732 5530 21788
rect 5530 21732 5534 21788
rect 5470 21728 5534 21732
rect 5550 21788 5614 21792
rect 5550 21732 5554 21788
rect 5554 21732 5610 21788
rect 5610 21732 5614 21788
rect 5550 21728 5614 21732
rect 5630 21788 5694 21792
rect 5630 21732 5634 21788
rect 5634 21732 5690 21788
rect 5690 21732 5694 21788
rect 5630 21728 5694 21732
rect 9829 21788 9893 21792
rect 9829 21732 9833 21788
rect 9833 21732 9889 21788
rect 9889 21732 9893 21788
rect 9829 21728 9893 21732
rect 9909 21788 9973 21792
rect 9909 21732 9913 21788
rect 9913 21732 9969 21788
rect 9969 21732 9973 21788
rect 9909 21728 9973 21732
rect 9989 21788 10053 21792
rect 9989 21732 9993 21788
rect 9993 21732 10049 21788
rect 10049 21732 10053 21788
rect 9989 21728 10053 21732
rect 10069 21788 10133 21792
rect 10069 21732 10073 21788
rect 10073 21732 10129 21788
rect 10129 21732 10133 21788
rect 10069 21728 10133 21732
rect 14268 21788 14332 21792
rect 14268 21732 14272 21788
rect 14272 21732 14328 21788
rect 14328 21732 14332 21788
rect 14268 21728 14332 21732
rect 14348 21788 14412 21792
rect 14348 21732 14352 21788
rect 14352 21732 14408 21788
rect 14408 21732 14412 21788
rect 14348 21728 14412 21732
rect 14428 21788 14492 21792
rect 14428 21732 14432 21788
rect 14432 21732 14488 21788
rect 14488 21732 14492 21788
rect 14428 21728 14492 21732
rect 14508 21788 14572 21792
rect 14508 21732 14512 21788
rect 14512 21732 14568 21788
rect 14568 21732 14572 21788
rect 14508 21728 14572 21732
rect 18707 21788 18771 21792
rect 18707 21732 18711 21788
rect 18711 21732 18767 21788
rect 18767 21732 18771 21788
rect 18707 21728 18771 21732
rect 18787 21788 18851 21792
rect 18787 21732 18791 21788
rect 18791 21732 18847 21788
rect 18847 21732 18851 21788
rect 18787 21728 18851 21732
rect 18867 21788 18931 21792
rect 18867 21732 18871 21788
rect 18871 21732 18927 21788
rect 18927 21732 18931 21788
rect 18867 21728 18931 21732
rect 18947 21788 19011 21792
rect 18947 21732 18951 21788
rect 18951 21732 19007 21788
rect 19007 21732 19011 21788
rect 18947 21728 19011 21732
rect 3171 21244 3235 21248
rect 3171 21188 3175 21244
rect 3175 21188 3231 21244
rect 3231 21188 3235 21244
rect 3171 21184 3235 21188
rect 3251 21244 3315 21248
rect 3251 21188 3255 21244
rect 3255 21188 3311 21244
rect 3311 21188 3315 21244
rect 3251 21184 3315 21188
rect 3331 21244 3395 21248
rect 3331 21188 3335 21244
rect 3335 21188 3391 21244
rect 3391 21188 3395 21244
rect 3331 21184 3395 21188
rect 3411 21244 3475 21248
rect 3411 21188 3415 21244
rect 3415 21188 3471 21244
rect 3471 21188 3475 21244
rect 3411 21184 3475 21188
rect 7610 21244 7674 21248
rect 7610 21188 7614 21244
rect 7614 21188 7670 21244
rect 7670 21188 7674 21244
rect 7610 21184 7674 21188
rect 7690 21244 7754 21248
rect 7690 21188 7694 21244
rect 7694 21188 7750 21244
rect 7750 21188 7754 21244
rect 7690 21184 7754 21188
rect 7770 21244 7834 21248
rect 7770 21188 7774 21244
rect 7774 21188 7830 21244
rect 7830 21188 7834 21244
rect 7770 21184 7834 21188
rect 7850 21244 7914 21248
rect 7850 21188 7854 21244
rect 7854 21188 7910 21244
rect 7910 21188 7914 21244
rect 7850 21184 7914 21188
rect 12049 21244 12113 21248
rect 12049 21188 12053 21244
rect 12053 21188 12109 21244
rect 12109 21188 12113 21244
rect 12049 21184 12113 21188
rect 12129 21244 12193 21248
rect 12129 21188 12133 21244
rect 12133 21188 12189 21244
rect 12189 21188 12193 21244
rect 12129 21184 12193 21188
rect 12209 21244 12273 21248
rect 12209 21188 12213 21244
rect 12213 21188 12269 21244
rect 12269 21188 12273 21244
rect 12209 21184 12273 21188
rect 12289 21244 12353 21248
rect 12289 21188 12293 21244
rect 12293 21188 12349 21244
rect 12349 21188 12353 21244
rect 12289 21184 12353 21188
rect 16488 21244 16552 21248
rect 16488 21188 16492 21244
rect 16492 21188 16548 21244
rect 16548 21188 16552 21244
rect 16488 21184 16552 21188
rect 16568 21244 16632 21248
rect 16568 21188 16572 21244
rect 16572 21188 16628 21244
rect 16628 21188 16632 21244
rect 16568 21184 16632 21188
rect 16648 21244 16712 21248
rect 16648 21188 16652 21244
rect 16652 21188 16708 21244
rect 16708 21188 16712 21244
rect 16648 21184 16712 21188
rect 16728 21244 16792 21248
rect 16728 21188 16732 21244
rect 16732 21188 16788 21244
rect 16788 21188 16792 21244
rect 16728 21184 16792 21188
rect 8156 20708 8220 20772
rect 5390 20700 5454 20704
rect 5390 20644 5394 20700
rect 5394 20644 5450 20700
rect 5450 20644 5454 20700
rect 5390 20640 5454 20644
rect 5470 20700 5534 20704
rect 5470 20644 5474 20700
rect 5474 20644 5530 20700
rect 5530 20644 5534 20700
rect 5470 20640 5534 20644
rect 5550 20700 5614 20704
rect 5550 20644 5554 20700
rect 5554 20644 5610 20700
rect 5610 20644 5614 20700
rect 5550 20640 5614 20644
rect 5630 20700 5694 20704
rect 5630 20644 5634 20700
rect 5634 20644 5690 20700
rect 5690 20644 5694 20700
rect 5630 20640 5694 20644
rect 9829 20700 9893 20704
rect 9829 20644 9833 20700
rect 9833 20644 9889 20700
rect 9889 20644 9893 20700
rect 9829 20640 9893 20644
rect 9909 20700 9973 20704
rect 9909 20644 9913 20700
rect 9913 20644 9969 20700
rect 9969 20644 9973 20700
rect 9909 20640 9973 20644
rect 9989 20700 10053 20704
rect 9989 20644 9993 20700
rect 9993 20644 10049 20700
rect 10049 20644 10053 20700
rect 9989 20640 10053 20644
rect 10069 20700 10133 20704
rect 10069 20644 10073 20700
rect 10073 20644 10129 20700
rect 10129 20644 10133 20700
rect 10069 20640 10133 20644
rect 14268 20700 14332 20704
rect 14268 20644 14272 20700
rect 14272 20644 14328 20700
rect 14328 20644 14332 20700
rect 14268 20640 14332 20644
rect 14348 20700 14412 20704
rect 14348 20644 14352 20700
rect 14352 20644 14408 20700
rect 14408 20644 14412 20700
rect 14348 20640 14412 20644
rect 14428 20700 14492 20704
rect 14428 20644 14432 20700
rect 14432 20644 14488 20700
rect 14488 20644 14492 20700
rect 14428 20640 14492 20644
rect 14508 20700 14572 20704
rect 14508 20644 14512 20700
rect 14512 20644 14568 20700
rect 14568 20644 14572 20700
rect 14508 20640 14572 20644
rect 18707 20700 18771 20704
rect 18707 20644 18711 20700
rect 18711 20644 18767 20700
rect 18767 20644 18771 20700
rect 18707 20640 18771 20644
rect 18787 20700 18851 20704
rect 18787 20644 18791 20700
rect 18791 20644 18847 20700
rect 18847 20644 18851 20700
rect 18787 20640 18851 20644
rect 18867 20700 18931 20704
rect 18867 20644 18871 20700
rect 18871 20644 18927 20700
rect 18927 20644 18931 20700
rect 18867 20640 18931 20644
rect 18947 20700 19011 20704
rect 18947 20644 18951 20700
rect 18951 20644 19007 20700
rect 19007 20644 19011 20700
rect 18947 20640 19011 20644
rect 3171 20156 3235 20160
rect 3171 20100 3175 20156
rect 3175 20100 3231 20156
rect 3231 20100 3235 20156
rect 3171 20096 3235 20100
rect 3251 20156 3315 20160
rect 3251 20100 3255 20156
rect 3255 20100 3311 20156
rect 3311 20100 3315 20156
rect 3251 20096 3315 20100
rect 3331 20156 3395 20160
rect 3331 20100 3335 20156
rect 3335 20100 3391 20156
rect 3391 20100 3395 20156
rect 3331 20096 3395 20100
rect 3411 20156 3475 20160
rect 3411 20100 3415 20156
rect 3415 20100 3471 20156
rect 3471 20100 3475 20156
rect 3411 20096 3475 20100
rect 7610 20156 7674 20160
rect 7610 20100 7614 20156
rect 7614 20100 7670 20156
rect 7670 20100 7674 20156
rect 7610 20096 7674 20100
rect 7690 20156 7754 20160
rect 7690 20100 7694 20156
rect 7694 20100 7750 20156
rect 7750 20100 7754 20156
rect 7690 20096 7754 20100
rect 7770 20156 7834 20160
rect 7770 20100 7774 20156
rect 7774 20100 7830 20156
rect 7830 20100 7834 20156
rect 7770 20096 7834 20100
rect 7850 20156 7914 20160
rect 7850 20100 7854 20156
rect 7854 20100 7910 20156
rect 7910 20100 7914 20156
rect 7850 20096 7914 20100
rect 12049 20156 12113 20160
rect 12049 20100 12053 20156
rect 12053 20100 12109 20156
rect 12109 20100 12113 20156
rect 12049 20096 12113 20100
rect 12129 20156 12193 20160
rect 12129 20100 12133 20156
rect 12133 20100 12189 20156
rect 12189 20100 12193 20156
rect 12129 20096 12193 20100
rect 12209 20156 12273 20160
rect 12209 20100 12213 20156
rect 12213 20100 12269 20156
rect 12269 20100 12273 20156
rect 12209 20096 12273 20100
rect 12289 20156 12353 20160
rect 12289 20100 12293 20156
rect 12293 20100 12349 20156
rect 12349 20100 12353 20156
rect 12289 20096 12353 20100
rect 16488 20156 16552 20160
rect 16488 20100 16492 20156
rect 16492 20100 16548 20156
rect 16548 20100 16552 20156
rect 16488 20096 16552 20100
rect 16568 20156 16632 20160
rect 16568 20100 16572 20156
rect 16572 20100 16628 20156
rect 16628 20100 16632 20156
rect 16568 20096 16632 20100
rect 16648 20156 16712 20160
rect 16648 20100 16652 20156
rect 16652 20100 16708 20156
rect 16708 20100 16712 20156
rect 16648 20096 16712 20100
rect 16728 20156 16792 20160
rect 16728 20100 16732 20156
rect 16732 20100 16788 20156
rect 16788 20100 16792 20156
rect 16728 20096 16792 20100
rect 5390 19612 5454 19616
rect 5390 19556 5394 19612
rect 5394 19556 5450 19612
rect 5450 19556 5454 19612
rect 5390 19552 5454 19556
rect 5470 19612 5534 19616
rect 5470 19556 5474 19612
rect 5474 19556 5530 19612
rect 5530 19556 5534 19612
rect 5470 19552 5534 19556
rect 5550 19612 5614 19616
rect 5550 19556 5554 19612
rect 5554 19556 5610 19612
rect 5610 19556 5614 19612
rect 5550 19552 5614 19556
rect 5630 19612 5694 19616
rect 5630 19556 5634 19612
rect 5634 19556 5690 19612
rect 5690 19556 5694 19612
rect 5630 19552 5694 19556
rect 9829 19612 9893 19616
rect 9829 19556 9833 19612
rect 9833 19556 9889 19612
rect 9889 19556 9893 19612
rect 9829 19552 9893 19556
rect 9909 19612 9973 19616
rect 9909 19556 9913 19612
rect 9913 19556 9969 19612
rect 9969 19556 9973 19612
rect 9909 19552 9973 19556
rect 9989 19612 10053 19616
rect 9989 19556 9993 19612
rect 9993 19556 10049 19612
rect 10049 19556 10053 19612
rect 9989 19552 10053 19556
rect 10069 19612 10133 19616
rect 10069 19556 10073 19612
rect 10073 19556 10129 19612
rect 10129 19556 10133 19612
rect 10069 19552 10133 19556
rect 14268 19612 14332 19616
rect 14268 19556 14272 19612
rect 14272 19556 14328 19612
rect 14328 19556 14332 19612
rect 14268 19552 14332 19556
rect 14348 19612 14412 19616
rect 14348 19556 14352 19612
rect 14352 19556 14408 19612
rect 14408 19556 14412 19612
rect 14348 19552 14412 19556
rect 14428 19612 14492 19616
rect 14428 19556 14432 19612
rect 14432 19556 14488 19612
rect 14488 19556 14492 19612
rect 14428 19552 14492 19556
rect 14508 19612 14572 19616
rect 14508 19556 14512 19612
rect 14512 19556 14568 19612
rect 14568 19556 14572 19612
rect 14508 19552 14572 19556
rect 18707 19612 18771 19616
rect 18707 19556 18711 19612
rect 18711 19556 18767 19612
rect 18767 19556 18771 19612
rect 18707 19552 18771 19556
rect 18787 19612 18851 19616
rect 18787 19556 18791 19612
rect 18791 19556 18847 19612
rect 18847 19556 18851 19612
rect 18787 19552 18851 19556
rect 18867 19612 18931 19616
rect 18867 19556 18871 19612
rect 18871 19556 18927 19612
rect 18927 19556 18931 19612
rect 18867 19552 18931 19556
rect 18947 19612 19011 19616
rect 18947 19556 18951 19612
rect 18951 19556 19007 19612
rect 19007 19556 19011 19612
rect 18947 19552 19011 19556
rect 2084 19408 2148 19412
rect 2084 19352 2098 19408
rect 2098 19352 2148 19408
rect 2084 19348 2148 19352
rect 3171 19068 3235 19072
rect 3171 19012 3175 19068
rect 3175 19012 3231 19068
rect 3231 19012 3235 19068
rect 3171 19008 3235 19012
rect 3251 19068 3315 19072
rect 3251 19012 3255 19068
rect 3255 19012 3311 19068
rect 3311 19012 3315 19068
rect 3251 19008 3315 19012
rect 3331 19068 3395 19072
rect 3331 19012 3335 19068
rect 3335 19012 3391 19068
rect 3391 19012 3395 19068
rect 3331 19008 3395 19012
rect 3411 19068 3475 19072
rect 3411 19012 3415 19068
rect 3415 19012 3471 19068
rect 3471 19012 3475 19068
rect 3411 19008 3475 19012
rect 7610 19068 7674 19072
rect 7610 19012 7614 19068
rect 7614 19012 7670 19068
rect 7670 19012 7674 19068
rect 7610 19008 7674 19012
rect 7690 19068 7754 19072
rect 7690 19012 7694 19068
rect 7694 19012 7750 19068
rect 7750 19012 7754 19068
rect 7690 19008 7754 19012
rect 7770 19068 7834 19072
rect 7770 19012 7774 19068
rect 7774 19012 7830 19068
rect 7830 19012 7834 19068
rect 7770 19008 7834 19012
rect 7850 19068 7914 19072
rect 7850 19012 7854 19068
rect 7854 19012 7910 19068
rect 7910 19012 7914 19068
rect 7850 19008 7914 19012
rect 12049 19068 12113 19072
rect 12049 19012 12053 19068
rect 12053 19012 12109 19068
rect 12109 19012 12113 19068
rect 12049 19008 12113 19012
rect 12129 19068 12193 19072
rect 12129 19012 12133 19068
rect 12133 19012 12189 19068
rect 12189 19012 12193 19068
rect 12129 19008 12193 19012
rect 12209 19068 12273 19072
rect 12209 19012 12213 19068
rect 12213 19012 12269 19068
rect 12269 19012 12273 19068
rect 12209 19008 12273 19012
rect 12289 19068 12353 19072
rect 12289 19012 12293 19068
rect 12293 19012 12349 19068
rect 12349 19012 12353 19068
rect 12289 19008 12353 19012
rect 16488 19068 16552 19072
rect 16488 19012 16492 19068
rect 16492 19012 16548 19068
rect 16548 19012 16552 19068
rect 16488 19008 16552 19012
rect 16568 19068 16632 19072
rect 16568 19012 16572 19068
rect 16572 19012 16628 19068
rect 16628 19012 16632 19068
rect 16568 19008 16632 19012
rect 16648 19068 16712 19072
rect 16648 19012 16652 19068
rect 16652 19012 16708 19068
rect 16708 19012 16712 19068
rect 16648 19008 16712 19012
rect 16728 19068 16792 19072
rect 16728 19012 16732 19068
rect 16732 19012 16788 19068
rect 16788 19012 16792 19068
rect 16728 19008 16792 19012
rect 5390 18524 5454 18528
rect 5390 18468 5394 18524
rect 5394 18468 5450 18524
rect 5450 18468 5454 18524
rect 5390 18464 5454 18468
rect 5470 18524 5534 18528
rect 5470 18468 5474 18524
rect 5474 18468 5530 18524
rect 5530 18468 5534 18524
rect 5470 18464 5534 18468
rect 5550 18524 5614 18528
rect 5550 18468 5554 18524
rect 5554 18468 5610 18524
rect 5610 18468 5614 18524
rect 5550 18464 5614 18468
rect 5630 18524 5694 18528
rect 5630 18468 5634 18524
rect 5634 18468 5690 18524
rect 5690 18468 5694 18524
rect 5630 18464 5694 18468
rect 9829 18524 9893 18528
rect 9829 18468 9833 18524
rect 9833 18468 9889 18524
rect 9889 18468 9893 18524
rect 9829 18464 9893 18468
rect 9909 18524 9973 18528
rect 9909 18468 9913 18524
rect 9913 18468 9969 18524
rect 9969 18468 9973 18524
rect 9909 18464 9973 18468
rect 9989 18524 10053 18528
rect 9989 18468 9993 18524
rect 9993 18468 10049 18524
rect 10049 18468 10053 18524
rect 9989 18464 10053 18468
rect 10069 18524 10133 18528
rect 10069 18468 10073 18524
rect 10073 18468 10129 18524
rect 10129 18468 10133 18524
rect 10069 18464 10133 18468
rect 14268 18524 14332 18528
rect 14268 18468 14272 18524
rect 14272 18468 14328 18524
rect 14328 18468 14332 18524
rect 14268 18464 14332 18468
rect 14348 18524 14412 18528
rect 14348 18468 14352 18524
rect 14352 18468 14408 18524
rect 14408 18468 14412 18524
rect 14348 18464 14412 18468
rect 14428 18524 14492 18528
rect 14428 18468 14432 18524
rect 14432 18468 14488 18524
rect 14488 18468 14492 18524
rect 14428 18464 14492 18468
rect 14508 18524 14572 18528
rect 14508 18468 14512 18524
rect 14512 18468 14568 18524
rect 14568 18468 14572 18524
rect 14508 18464 14572 18468
rect 18707 18524 18771 18528
rect 18707 18468 18711 18524
rect 18711 18468 18767 18524
rect 18767 18468 18771 18524
rect 18707 18464 18771 18468
rect 18787 18524 18851 18528
rect 18787 18468 18791 18524
rect 18791 18468 18847 18524
rect 18847 18468 18851 18524
rect 18787 18464 18851 18468
rect 18867 18524 18931 18528
rect 18867 18468 18871 18524
rect 18871 18468 18927 18524
rect 18927 18468 18931 18524
rect 18867 18464 18931 18468
rect 18947 18524 19011 18528
rect 18947 18468 18951 18524
rect 18951 18468 19007 18524
rect 19007 18468 19011 18524
rect 18947 18464 19011 18468
rect 3171 17980 3235 17984
rect 3171 17924 3175 17980
rect 3175 17924 3231 17980
rect 3231 17924 3235 17980
rect 3171 17920 3235 17924
rect 3251 17980 3315 17984
rect 3251 17924 3255 17980
rect 3255 17924 3311 17980
rect 3311 17924 3315 17980
rect 3251 17920 3315 17924
rect 3331 17980 3395 17984
rect 3331 17924 3335 17980
rect 3335 17924 3391 17980
rect 3391 17924 3395 17980
rect 3331 17920 3395 17924
rect 3411 17980 3475 17984
rect 3411 17924 3415 17980
rect 3415 17924 3471 17980
rect 3471 17924 3475 17980
rect 3411 17920 3475 17924
rect 7610 17980 7674 17984
rect 7610 17924 7614 17980
rect 7614 17924 7670 17980
rect 7670 17924 7674 17980
rect 7610 17920 7674 17924
rect 7690 17980 7754 17984
rect 7690 17924 7694 17980
rect 7694 17924 7750 17980
rect 7750 17924 7754 17980
rect 7690 17920 7754 17924
rect 7770 17980 7834 17984
rect 7770 17924 7774 17980
rect 7774 17924 7830 17980
rect 7830 17924 7834 17980
rect 7770 17920 7834 17924
rect 7850 17980 7914 17984
rect 7850 17924 7854 17980
rect 7854 17924 7910 17980
rect 7910 17924 7914 17980
rect 7850 17920 7914 17924
rect 12049 17980 12113 17984
rect 12049 17924 12053 17980
rect 12053 17924 12109 17980
rect 12109 17924 12113 17980
rect 12049 17920 12113 17924
rect 12129 17980 12193 17984
rect 12129 17924 12133 17980
rect 12133 17924 12189 17980
rect 12189 17924 12193 17980
rect 12129 17920 12193 17924
rect 12209 17980 12273 17984
rect 12209 17924 12213 17980
rect 12213 17924 12269 17980
rect 12269 17924 12273 17980
rect 12209 17920 12273 17924
rect 12289 17980 12353 17984
rect 12289 17924 12293 17980
rect 12293 17924 12349 17980
rect 12349 17924 12353 17980
rect 12289 17920 12353 17924
rect 16488 17980 16552 17984
rect 16488 17924 16492 17980
rect 16492 17924 16548 17980
rect 16548 17924 16552 17980
rect 16488 17920 16552 17924
rect 16568 17980 16632 17984
rect 16568 17924 16572 17980
rect 16572 17924 16628 17980
rect 16628 17924 16632 17980
rect 16568 17920 16632 17924
rect 16648 17980 16712 17984
rect 16648 17924 16652 17980
rect 16652 17924 16708 17980
rect 16708 17924 16712 17980
rect 16648 17920 16712 17924
rect 16728 17980 16792 17984
rect 16728 17924 16732 17980
rect 16732 17924 16788 17980
rect 16788 17924 16792 17980
rect 16728 17920 16792 17924
rect 5390 17436 5454 17440
rect 5390 17380 5394 17436
rect 5394 17380 5450 17436
rect 5450 17380 5454 17436
rect 5390 17376 5454 17380
rect 5470 17436 5534 17440
rect 5470 17380 5474 17436
rect 5474 17380 5530 17436
rect 5530 17380 5534 17436
rect 5470 17376 5534 17380
rect 5550 17436 5614 17440
rect 5550 17380 5554 17436
rect 5554 17380 5610 17436
rect 5610 17380 5614 17436
rect 5550 17376 5614 17380
rect 5630 17436 5694 17440
rect 5630 17380 5634 17436
rect 5634 17380 5690 17436
rect 5690 17380 5694 17436
rect 5630 17376 5694 17380
rect 9829 17436 9893 17440
rect 9829 17380 9833 17436
rect 9833 17380 9889 17436
rect 9889 17380 9893 17436
rect 9829 17376 9893 17380
rect 9909 17436 9973 17440
rect 9909 17380 9913 17436
rect 9913 17380 9969 17436
rect 9969 17380 9973 17436
rect 9909 17376 9973 17380
rect 9989 17436 10053 17440
rect 9989 17380 9993 17436
rect 9993 17380 10049 17436
rect 10049 17380 10053 17436
rect 9989 17376 10053 17380
rect 10069 17436 10133 17440
rect 10069 17380 10073 17436
rect 10073 17380 10129 17436
rect 10129 17380 10133 17436
rect 10069 17376 10133 17380
rect 14268 17436 14332 17440
rect 14268 17380 14272 17436
rect 14272 17380 14328 17436
rect 14328 17380 14332 17436
rect 14268 17376 14332 17380
rect 14348 17436 14412 17440
rect 14348 17380 14352 17436
rect 14352 17380 14408 17436
rect 14408 17380 14412 17436
rect 14348 17376 14412 17380
rect 14428 17436 14492 17440
rect 14428 17380 14432 17436
rect 14432 17380 14488 17436
rect 14488 17380 14492 17436
rect 14428 17376 14492 17380
rect 14508 17436 14572 17440
rect 14508 17380 14512 17436
rect 14512 17380 14568 17436
rect 14568 17380 14572 17436
rect 14508 17376 14572 17380
rect 18707 17436 18771 17440
rect 18707 17380 18711 17436
rect 18711 17380 18767 17436
rect 18767 17380 18771 17436
rect 18707 17376 18771 17380
rect 18787 17436 18851 17440
rect 18787 17380 18791 17436
rect 18791 17380 18847 17436
rect 18847 17380 18851 17436
rect 18787 17376 18851 17380
rect 18867 17436 18931 17440
rect 18867 17380 18871 17436
rect 18871 17380 18927 17436
rect 18927 17380 18931 17436
rect 18867 17376 18931 17380
rect 18947 17436 19011 17440
rect 18947 17380 18951 17436
rect 18951 17380 19007 17436
rect 19007 17380 19011 17436
rect 18947 17376 19011 17380
rect 3924 17232 3988 17236
rect 3924 17176 3974 17232
rect 3974 17176 3988 17232
rect 3924 17172 3988 17176
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 3004 16628 3068 16692
rect 5390 16348 5454 16352
rect 5390 16292 5394 16348
rect 5394 16292 5450 16348
rect 5450 16292 5454 16348
rect 5390 16288 5454 16292
rect 5470 16348 5534 16352
rect 5470 16292 5474 16348
rect 5474 16292 5530 16348
rect 5530 16292 5534 16348
rect 5470 16288 5534 16292
rect 5550 16348 5614 16352
rect 5550 16292 5554 16348
rect 5554 16292 5610 16348
rect 5610 16292 5614 16348
rect 5550 16288 5614 16292
rect 5630 16348 5694 16352
rect 5630 16292 5634 16348
rect 5634 16292 5690 16348
rect 5690 16292 5694 16348
rect 5630 16288 5694 16292
rect 9829 16348 9893 16352
rect 9829 16292 9833 16348
rect 9833 16292 9889 16348
rect 9889 16292 9893 16348
rect 9829 16288 9893 16292
rect 9909 16348 9973 16352
rect 9909 16292 9913 16348
rect 9913 16292 9969 16348
rect 9969 16292 9973 16348
rect 9909 16288 9973 16292
rect 9989 16348 10053 16352
rect 9989 16292 9993 16348
rect 9993 16292 10049 16348
rect 10049 16292 10053 16348
rect 9989 16288 10053 16292
rect 10069 16348 10133 16352
rect 10069 16292 10073 16348
rect 10073 16292 10129 16348
rect 10129 16292 10133 16348
rect 10069 16288 10133 16292
rect 14268 16348 14332 16352
rect 14268 16292 14272 16348
rect 14272 16292 14328 16348
rect 14328 16292 14332 16348
rect 14268 16288 14332 16292
rect 14348 16348 14412 16352
rect 14348 16292 14352 16348
rect 14352 16292 14408 16348
rect 14408 16292 14412 16348
rect 14348 16288 14412 16292
rect 14428 16348 14492 16352
rect 14428 16292 14432 16348
rect 14432 16292 14488 16348
rect 14488 16292 14492 16348
rect 14428 16288 14492 16292
rect 14508 16348 14572 16352
rect 14508 16292 14512 16348
rect 14512 16292 14568 16348
rect 14568 16292 14572 16348
rect 14508 16288 14572 16292
rect 18707 16348 18771 16352
rect 18707 16292 18711 16348
rect 18711 16292 18767 16348
rect 18767 16292 18771 16348
rect 18707 16288 18771 16292
rect 18787 16348 18851 16352
rect 18787 16292 18791 16348
rect 18791 16292 18847 16348
rect 18847 16292 18851 16348
rect 18787 16288 18851 16292
rect 18867 16348 18931 16352
rect 18867 16292 18871 16348
rect 18871 16292 18927 16348
rect 18927 16292 18931 16348
rect 18867 16288 18931 16292
rect 18947 16348 19011 16352
rect 18947 16292 18951 16348
rect 18951 16292 19007 16348
rect 19007 16292 19011 16348
rect 18947 16288 19011 16292
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 5390 15260 5454 15264
rect 5390 15204 5394 15260
rect 5394 15204 5450 15260
rect 5450 15204 5454 15260
rect 5390 15200 5454 15204
rect 5470 15260 5534 15264
rect 5470 15204 5474 15260
rect 5474 15204 5530 15260
rect 5530 15204 5534 15260
rect 5470 15200 5534 15204
rect 5550 15260 5614 15264
rect 5550 15204 5554 15260
rect 5554 15204 5610 15260
rect 5610 15204 5614 15260
rect 5550 15200 5614 15204
rect 5630 15260 5694 15264
rect 5630 15204 5634 15260
rect 5634 15204 5690 15260
rect 5690 15204 5694 15260
rect 5630 15200 5694 15204
rect 9829 15260 9893 15264
rect 9829 15204 9833 15260
rect 9833 15204 9889 15260
rect 9889 15204 9893 15260
rect 9829 15200 9893 15204
rect 9909 15260 9973 15264
rect 9909 15204 9913 15260
rect 9913 15204 9969 15260
rect 9969 15204 9973 15260
rect 9909 15200 9973 15204
rect 9989 15260 10053 15264
rect 9989 15204 9993 15260
rect 9993 15204 10049 15260
rect 10049 15204 10053 15260
rect 9989 15200 10053 15204
rect 10069 15260 10133 15264
rect 10069 15204 10073 15260
rect 10073 15204 10129 15260
rect 10129 15204 10133 15260
rect 10069 15200 10133 15204
rect 14268 15260 14332 15264
rect 14268 15204 14272 15260
rect 14272 15204 14328 15260
rect 14328 15204 14332 15260
rect 14268 15200 14332 15204
rect 14348 15260 14412 15264
rect 14348 15204 14352 15260
rect 14352 15204 14408 15260
rect 14408 15204 14412 15260
rect 14348 15200 14412 15204
rect 14428 15260 14492 15264
rect 14428 15204 14432 15260
rect 14432 15204 14488 15260
rect 14488 15204 14492 15260
rect 14428 15200 14492 15204
rect 14508 15260 14572 15264
rect 14508 15204 14512 15260
rect 14512 15204 14568 15260
rect 14568 15204 14572 15260
rect 14508 15200 14572 15204
rect 18707 15260 18771 15264
rect 18707 15204 18711 15260
rect 18711 15204 18767 15260
rect 18767 15204 18771 15260
rect 18707 15200 18771 15204
rect 18787 15260 18851 15264
rect 18787 15204 18791 15260
rect 18791 15204 18847 15260
rect 18847 15204 18851 15260
rect 18787 15200 18851 15204
rect 18867 15260 18931 15264
rect 18867 15204 18871 15260
rect 18871 15204 18927 15260
rect 18927 15204 18931 15260
rect 18867 15200 18931 15204
rect 18947 15260 19011 15264
rect 18947 15204 18951 15260
rect 18951 15204 19007 15260
rect 19007 15204 19011 15260
rect 18947 15200 19011 15204
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 5390 14172 5454 14176
rect 5390 14116 5394 14172
rect 5394 14116 5450 14172
rect 5450 14116 5454 14172
rect 5390 14112 5454 14116
rect 5470 14172 5534 14176
rect 5470 14116 5474 14172
rect 5474 14116 5530 14172
rect 5530 14116 5534 14172
rect 5470 14112 5534 14116
rect 5550 14172 5614 14176
rect 5550 14116 5554 14172
rect 5554 14116 5610 14172
rect 5610 14116 5614 14172
rect 5550 14112 5614 14116
rect 5630 14172 5694 14176
rect 5630 14116 5634 14172
rect 5634 14116 5690 14172
rect 5690 14116 5694 14172
rect 5630 14112 5694 14116
rect 9829 14172 9893 14176
rect 9829 14116 9833 14172
rect 9833 14116 9889 14172
rect 9889 14116 9893 14172
rect 9829 14112 9893 14116
rect 9909 14172 9973 14176
rect 9909 14116 9913 14172
rect 9913 14116 9969 14172
rect 9969 14116 9973 14172
rect 9909 14112 9973 14116
rect 9989 14172 10053 14176
rect 9989 14116 9993 14172
rect 9993 14116 10049 14172
rect 10049 14116 10053 14172
rect 9989 14112 10053 14116
rect 10069 14172 10133 14176
rect 10069 14116 10073 14172
rect 10073 14116 10129 14172
rect 10129 14116 10133 14172
rect 10069 14112 10133 14116
rect 14268 14172 14332 14176
rect 14268 14116 14272 14172
rect 14272 14116 14328 14172
rect 14328 14116 14332 14172
rect 14268 14112 14332 14116
rect 14348 14172 14412 14176
rect 14348 14116 14352 14172
rect 14352 14116 14408 14172
rect 14408 14116 14412 14172
rect 14348 14112 14412 14116
rect 14428 14172 14492 14176
rect 14428 14116 14432 14172
rect 14432 14116 14488 14172
rect 14488 14116 14492 14172
rect 14428 14112 14492 14116
rect 14508 14172 14572 14176
rect 14508 14116 14512 14172
rect 14512 14116 14568 14172
rect 14568 14116 14572 14172
rect 14508 14112 14572 14116
rect 18707 14172 18771 14176
rect 18707 14116 18711 14172
rect 18711 14116 18767 14172
rect 18767 14116 18771 14172
rect 18707 14112 18771 14116
rect 18787 14172 18851 14176
rect 18787 14116 18791 14172
rect 18791 14116 18847 14172
rect 18847 14116 18851 14172
rect 18787 14112 18851 14116
rect 18867 14172 18931 14176
rect 18867 14116 18871 14172
rect 18871 14116 18927 14172
rect 18927 14116 18931 14172
rect 18867 14112 18931 14116
rect 18947 14172 19011 14176
rect 18947 14116 18951 14172
rect 18951 14116 19007 14172
rect 19007 14116 19011 14172
rect 18947 14112 19011 14116
rect 2084 13772 2148 13836
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 5390 13084 5454 13088
rect 5390 13028 5394 13084
rect 5394 13028 5450 13084
rect 5450 13028 5454 13084
rect 5390 13024 5454 13028
rect 5470 13084 5534 13088
rect 5470 13028 5474 13084
rect 5474 13028 5530 13084
rect 5530 13028 5534 13084
rect 5470 13024 5534 13028
rect 5550 13084 5614 13088
rect 5550 13028 5554 13084
rect 5554 13028 5610 13084
rect 5610 13028 5614 13084
rect 5550 13024 5614 13028
rect 5630 13084 5694 13088
rect 5630 13028 5634 13084
rect 5634 13028 5690 13084
rect 5690 13028 5694 13084
rect 5630 13024 5694 13028
rect 9829 13084 9893 13088
rect 9829 13028 9833 13084
rect 9833 13028 9889 13084
rect 9889 13028 9893 13084
rect 9829 13024 9893 13028
rect 9909 13084 9973 13088
rect 9909 13028 9913 13084
rect 9913 13028 9969 13084
rect 9969 13028 9973 13084
rect 9909 13024 9973 13028
rect 9989 13084 10053 13088
rect 9989 13028 9993 13084
rect 9993 13028 10049 13084
rect 10049 13028 10053 13084
rect 9989 13024 10053 13028
rect 10069 13084 10133 13088
rect 10069 13028 10073 13084
rect 10073 13028 10129 13084
rect 10129 13028 10133 13084
rect 10069 13024 10133 13028
rect 14268 13084 14332 13088
rect 14268 13028 14272 13084
rect 14272 13028 14328 13084
rect 14328 13028 14332 13084
rect 14268 13024 14332 13028
rect 14348 13084 14412 13088
rect 14348 13028 14352 13084
rect 14352 13028 14408 13084
rect 14408 13028 14412 13084
rect 14348 13024 14412 13028
rect 14428 13084 14492 13088
rect 14428 13028 14432 13084
rect 14432 13028 14488 13084
rect 14488 13028 14492 13084
rect 14428 13024 14492 13028
rect 14508 13084 14572 13088
rect 14508 13028 14512 13084
rect 14512 13028 14568 13084
rect 14568 13028 14572 13084
rect 14508 13024 14572 13028
rect 18707 13084 18771 13088
rect 18707 13028 18711 13084
rect 18711 13028 18767 13084
rect 18767 13028 18771 13084
rect 18707 13024 18771 13028
rect 18787 13084 18851 13088
rect 18787 13028 18791 13084
rect 18791 13028 18847 13084
rect 18847 13028 18851 13084
rect 18787 13024 18851 13028
rect 18867 13084 18931 13088
rect 18867 13028 18871 13084
rect 18871 13028 18927 13084
rect 18927 13028 18931 13084
rect 18867 13024 18931 13028
rect 18947 13084 19011 13088
rect 18947 13028 18951 13084
rect 18951 13028 19007 13084
rect 19007 13028 19011 13084
rect 18947 13024 19011 13028
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 5390 11996 5454 12000
rect 5390 11940 5394 11996
rect 5394 11940 5450 11996
rect 5450 11940 5454 11996
rect 5390 11936 5454 11940
rect 5470 11996 5534 12000
rect 5470 11940 5474 11996
rect 5474 11940 5530 11996
rect 5530 11940 5534 11996
rect 5470 11936 5534 11940
rect 5550 11996 5614 12000
rect 5550 11940 5554 11996
rect 5554 11940 5610 11996
rect 5610 11940 5614 11996
rect 5550 11936 5614 11940
rect 5630 11996 5694 12000
rect 5630 11940 5634 11996
rect 5634 11940 5690 11996
rect 5690 11940 5694 11996
rect 5630 11936 5694 11940
rect 9829 11996 9893 12000
rect 9829 11940 9833 11996
rect 9833 11940 9889 11996
rect 9889 11940 9893 11996
rect 9829 11936 9893 11940
rect 9909 11996 9973 12000
rect 9909 11940 9913 11996
rect 9913 11940 9969 11996
rect 9969 11940 9973 11996
rect 9909 11936 9973 11940
rect 9989 11996 10053 12000
rect 9989 11940 9993 11996
rect 9993 11940 10049 11996
rect 10049 11940 10053 11996
rect 9989 11936 10053 11940
rect 10069 11996 10133 12000
rect 10069 11940 10073 11996
rect 10073 11940 10129 11996
rect 10129 11940 10133 11996
rect 10069 11936 10133 11940
rect 14268 11996 14332 12000
rect 14268 11940 14272 11996
rect 14272 11940 14328 11996
rect 14328 11940 14332 11996
rect 14268 11936 14332 11940
rect 14348 11996 14412 12000
rect 14348 11940 14352 11996
rect 14352 11940 14408 11996
rect 14408 11940 14412 11996
rect 14348 11936 14412 11940
rect 14428 11996 14492 12000
rect 14428 11940 14432 11996
rect 14432 11940 14488 11996
rect 14488 11940 14492 11996
rect 14428 11936 14492 11940
rect 14508 11996 14572 12000
rect 14508 11940 14512 11996
rect 14512 11940 14568 11996
rect 14568 11940 14572 11996
rect 14508 11936 14572 11940
rect 18707 11996 18771 12000
rect 18707 11940 18711 11996
rect 18711 11940 18767 11996
rect 18767 11940 18771 11996
rect 18707 11936 18771 11940
rect 18787 11996 18851 12000
rect 18787 11940 18791 11996
rect 18791 11940 18847 11996
rect 18847 11940 18851 11996
rect 18787 11936 18851 11940
rect 18867 11996 18931 12000
rect 18867 11940 18871 11996
rect 18871 11940 18927 11996
rect 18927 11940 18931 11996
rect 18867 11936 18931 11940
rect 18947 11996 19011 12000
rect 18947 11940 18951 11996
rect 18951 11940 19007 11996
rect 19007 11940 19011 11996
rect 18947 11936 19011 11940
rect 1900 11596 1964 11660
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 4292 10976 4356 10980
rect 4292 10920 4306 10976
rect 4306 10920 4356 10976
rect 4292 10916 4356 10920
rect 5390 10908 5454 10912
rect 5390 10852 5394 10908
rect 5394 10852 5450 10908
rect 5450 10852 5454 10908
rect 5390 10848 5454 10852
rect 5470 10908 5534 10912
rect 5470 10852 5474 10908
rect 5474 10852 5530 10908
rect 5530 10852 5534 10908
rect 5470 10848 5534 10852
rect 5550 10908 5614 10912
rect 5550 10852 5554 10908
rect 5554 10852 5610 10908
rect 5610 10852 5614 10908
rect 5550 10848 5614 10852
rect 5630 10908 5694 10912
rect 5630 10852 5634 10908
rect 5634 10852 5690 10908
rect 5690 10852 5694 10908
rect 5630 10848 5694 10852
rect 9829 10908 9893 10912
rect 9829 10852 9833 10908
rect 9833 10852 9889 10908
rect 9889 10852 9893 10908
rect 9829 10848 9893 10852
rect 9909 10908 9973 10912
rect 9909 10852 9913 10908
rect 9913 10852 9969 10908
rect 9969 10852 9973 10908
rect 9909 10848 9973 10852
rect 9989 10908 10053 10912
rect 9989 10852 9993 10908
rect 9993 10852 10049 10908
rect 10049 10852 10053 10908
rect 9989 10848 10053 10852
rect 10069 10908 10133 10912
rect 10069 10852 10073 10908
rect 10073 10852 10129 10908
rect 10129 10852 10133 10908
rect 10069 10848 10133 10852
rect 14268 10908 14332 10912
rect 14268 10852 14272 10908
rect 14272 10852 14328 10908
rect 14328 10852 14332 10908
rect 14268 10848 14332 10852
rect 14348 10908 14412 10912
rect 14348 10852 14352 10908
rect 14352 10852 14408 10908
rect 14408 10852 14412 10908
rect 14348 10848 14412 10852
rect 14428 10908 14492 10912
rect 14428 10852 14432 10908
rect 14432 10852 14488 10908
rect 14488 10852 14492 10908
rect 14428 10848 14492 10852
rect 14508 10908 14572 10912
rect 14508 10852 14512 10908
rect 14512 10852 14568 10908
rect 14568 10852 14572 10908
rect 14508 10848 14572 10852
rect 18707 10908 18771 10912
rect 18707 10852 18711 10908
rect 18711 10852 18767 10908
rect 18767 10852 18771 10908
rect 18707 10848 18771 10852
rect 18787 10908 18851 10912
rect 18787 10852 18791 10908
rect 18791 10852 18847 10908
rect 18847 10852 18851 10908
rect 18787 10848 18851 10852
rect 18867 10908 18931 10912
rect 18867 10852 18871 10908
rect 18871 10852 18927 10908
rect 18927 10852 18931 10908
rect 18867 10848 18931 10852
rect 18947 10908 19011 10912
rect 18947 10852 18951 10908
rect 18951 10852 19007 10908
rect 19007 10852 19011 10908
rect 18947 10848 19011 10852
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 5390 9820 5454 9824
rect 5390 9764 5394 9820
rect 5394 9764 5450 9820
rect 5450 9764 5454 9820
rect 5390 9760 5454 9764
rect 5470 9820 5534 9824
rect 5470 9764 5474 9820
rect 5474 9764 5530 9820
rect 5530 9764 5534 9820
rect 5470 9760 5534 9764
rect 5550 9820 5614 9824
rect 5550 9764 5554 9820
rect 5554 9764 5610 9820
rect 5610 9764 5614 9820
rect 5550 9760 5614 9764
rect 5630 9820 5694 9824
rect 5630 9764 5634 9820
rect 5634 9764 5690 9820
rect 5690 9764 5694 9820
rect 5630 9760 5694 9764
rect 9829 9820 9893 9824
rect 9829 9764 9833 9820
rect 9833 9764 9889 9820
rect 9889 9764 9893 9820
rect 9829 9760 9893 9764
rect 9909 9820 9973 9824
rect 9909 9764 9913 9820
rect 9913 9764 9969 9820
rect 9969 9764 9973 9820
rect 9909 9760 9973 9764
rect 9989 9820 10053 9824
rect 9989 9764 9993 9820
rect 9993 9764 10049 9820
rect 10049 9764 10053 9820
rect 9989 9760 10053 9764
rect 10069 9820 10133 9824
rect 10069 9764 10073 9820
rect 10073 9764 10129 9820
rect 10129 9764 10133 9820
rect 10069 9760 10133 9764
rect 14268 9820 14332 9824
rect 14268 9764 14272 9820
rect 14272 9764 14328 9820
rect 14328 9764 14332 9820
rect 14268 9760 14332 9764
rect 14348 9820 14412 9824
rect 14348 9764 14352 9820
rect 14352 9764 14408 9820
rect 14408 9764 14412 9820
rect 14348 9760 14412 9764
rect 14428 9820 14492 9824
rect 14428 9764 14432 9820
rect 14432 9764 14488 9820
rect 14488 9764 14492 9820
rect 14428 9760 14492 9764
rect 14508 9820 14572 9824
rect 14508 9764 14512 9820
rect 14512 9764 14568 9820
rect 14568 9764 14572 9820
rect 14508 9760 14572 9764
rect 18707 9820 18771 9824
rect 18707 9764 18711 9820
rect 18711 9764 18767 9820
rect 18767 9764 18771 9820
rect 18707 9760 18771 9764
rect 18787 9820 18851 9824
rect 18787 9764 18791 9820
rect 18791 9764 18847 9820
rect 18847 9764 18851 9820
rect 18787 9760 18851 9764
rect 18867 9820 18931 9824
rect 18867 9764 18871 9820
rect 18871 9764 18927 9820
rect 18927 9764 18931 9820
rect 18867 9760 18931 9764
rect 18947 9820 19011 9824
rect 18947 9764 18951 9820
rect 18951 9764 19007 9820
rect 19007 9764 19011 9820
rect 18947 9760 19011 9764
rect 3004 9692 3068 9756
rect 4660 9556 4724 9620
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 5390 8732 5454 8736
rect 5390 8676 5394 8732
rect 5394 8676 5450 8732
rect 5450 8676 5454 8732
rect 5390 8672 5454 8676
rect 5470 8732 5534 8736
rect 5470 8676 5474 8732
rect 5474 8676 5530 8732
rect 5530 8676 5534 8732
rect 5470 8672 5534 8676
rect 5550 8732 5614 8736
rect 5550 8676 5554 8732
rect 5554 8676 5610 8732
rect 5610 8676 5614 8732
rect 5550 8672 5614 8676
rect 5630 8732 5694 8736
rect 5630 8676 5634 8732
rect 5634 8676 5690 8732
rect 5690 8676 5694 8732
rect 5630 8672 5694 8676
rect 9829 8732 9893 8736
rect 9829 8676 9833 8732
rect 9833 8676 9889 8732
rect 9889 8676 9893 8732
rect 9829 8672 9893 8676
rect 9909 8732 9973 8736
rect 9909 8676 9913 8732
rect 9913 8676 9969 8732
rect 9969 8676 9973 8732
rect 9909 8672 9973 8676
rect 9989 8732 10053 8736
rect 9989 8676 9993 8732
rect 9993 8676 10049 8732
rect 10049 8676 10053 8732
rect 9989 8672 10053 8676
rect 10069 8732 10133 8736
rect 10069 8676 10073 8732
rect 10073 8676 10129 8732
rect 10129 8676 10133 8732
rect 10069 8672 10133 8676
rect 14268 8732 14332 8736
rect 14268 8676 14272 8732
rect 14272 8676 14328 8732
rect 14328 8676 14332 8732
rect 14268 8672 14332 8676
rect 14348 8732 14412 8736
rect 14348 8676 14352 8732
rect 14352 8676 14408 8732
rect 14408 8676 14412 8732
rect 14348 8672 14412 8676
rect 14428 8732 14492 8736
rect 14428 8676 14432 8732
rect 14432 8676 14488 8732
rect 14488 8676 14492 8732
rect 14428 8672 14492 8676
rect 14508 8732 14572 8736
rect 14508 8676 14512 8732
rect 14512 8676 14568 8732
rect 14568 8676 14572 8732
rect 14508 8672 14572 8676
rect 18707 8732 18771 8736
rect 18707 8676 18711 8732
rect 18711 8676 18767 8732
rect 18767 8676 18771 8732
rect 18707 8672 18771 8676
rect 18787 8732 18851 8736
rect 18787 8676 18791 8732
rect 18791 8676 18847 8732
rect 18847 8676 18851 8732
rect 18787 8672 18851 8676
rect 18867 8732 18931 8736
rect 18867 8676 18871 8732
rect 18871 8676 18927 8732
rect 18927 8676 18931 8732
rect 18867 8672 18931 8676
rect 18947 8732 19011 8736
rect 18947 8676 18951 8732
rect 18951 8676 19007 8732
rect 19007 8676 19011 8732
rect 18947 8672 19011 8676
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 6684 6564 6748 6628
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 4844 5536 4908 5540
rect 4844 5480 4858 5536
rect 4858 5480 4908 5536
rect 4844 5476 4908 5480
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 3163 47360 3483 47376
rect 3163 47296 3171 47360
rect 3235 47296 3251 47360
rect 3315 47296 3331 47360
rect 3395 47296 3411 47360
rect 3475 47296 3483 47360
rect 3163 46272 3483 47296
rect 3163 46208 3171 46272
rect 3235 46208 3251 46272
rect 3315 46208 3331 46272
rect 3395 46208 3411 46272
rect 3475 46208 3483 46272
rect 3163 45184 3483 46208
rect 3163 45120 3171 45184
rect 3235 45120 3251 45184
rect 3315 45120 3331 45184
rect 3395 45120 3411 45184
rect 3475 45120 3483 45184
rect 3163 44096 3483 45120
rect 3163 44032 3171 44096
rect 3235 44032 3251 44096
rect 3315 44032 3331 44096
rect 3395 44032 3411 44096
rect 3475 44032 3483 44096
rect 3163 43008 3483 44032
rect 3163 42944 3171 43008
rect 3235 42944 3251 43008
rect 3315 42944 3331 43008
rect 3395 42944 3411 43008
rect 3475 42944 3483 43008
rect 3163 41920 3483 42944
rect 3163 41856 3171 41920
rect 3235 41856 3251 41920
rect 3315 41856 3331 41920
rect 3395 41856 3411 41920
rect 3475 41856 3483 41920
rect 3163 40832 3483 41856
rect 3163 40768 3171 40832
rect 3235 40768 3251 40832
rect 3315 40768 3331 40832
rect 3395 40768 3411 40832
rect 3475 40768 3483 40832
rect 3163 39744 3483 40768
rect 3163 39680 3171 39744
rect 3235 39680 3251 39744
rect 3315 39680 3331 39744
rect 3395 39680 3411 39744
rect 3475 39680 3483 39744
rect 3163 38656 3483 39680
rect 3163 38592 3171 38656
rect 3235 38592 3251 38656
rect 3315 38592 3331 38656
rect 3395 38592 3411 38656
rect 3475 38592 3483 38656
rect 3163 37568 3483 38592
rect 3163 37504 3171 37568
rect 3235 37504 3251 37568
rect 3315 37504 3331 37568
rect 3395 37504 3411 37568
rect 3475 37504 3483 37568
rect 3163 36480 3483 37504
rect 3163 36416 3171 36480
rect 3235 36416 3251 36480
rect 3315 36416 3331 36480
rect 3395 36416 3411 36480
rect 3475 36416 3483 36480
rect 3163 35392 3483 36416
rect 3163 35328 3171 35392
rect 3235 35328 3251 35392
rect 3315 35328 3331 35392
rect 3395 35328 3411 35392
rect 3475 35328 3483 35392
rect 3163 34304 3483 35328
rect 3163 34240 3171 34304
rect 3235 34240 3251 34304
rect 3315 34240 3331 34304
rect 3395 34240 3411 34304
rect 3475 34240 3483 34304
rect 3163 33216 3483 34240
rect 3163 33152 3171 33216
rect 3235 33152 3251 33216
rect 3315 33152 3331 33216
rect 3395 33152 3411 33216
rect 3475 33152 3483 33216
rect 3163 32128 3483 33152
rect 3163 32064 3171 32128
rect 3235 32064 3251 32128
rect 3315 32064 3331 32128
rect 3395 32064 3411 32128
rect 3475 32064 3483 32128
rect 3163 31040 3483 32064
rect 3163 30976 3171 31040
rect 3235 30976 3251 31040
rect 3315 30976 3331 31040
rect 3395 30976 3411 31040
rect 3475 30976 3483 31040
rect 3163 29952 3483 30976
rect 5382 46816 5702 47376
rect 5382 46752 5390 46816
rect 5454 46752 5470 46816
rect 5534 46752 5550 46816
rect 5614 46752 5630 46816
rect 5694 46752 5702 46816
rect 5382 45728 5702 46752
rect 5382 45664 5390 45728
rect 5454 45664 5470 45728
rect 5534 45664 5550 45728
rect 5614 45664 5630 45728
rect 5694 45664 5702 45728
rect 5382 44640 5702 45664
rect 5382 44576 5390 44640
rect 5454 44576 5470 44640
rect 5534 44576 5550 44640
rect 5614 44576 5630 44640
rect 5694 44576 5702 44640
rect 5382 43552 5702 44576
rect 5382 43488 5390 43552
rect 5454 43488 5470 43552
rect 5534 43488 5550 43552
rect 5614 43488 5630 43552
rect 5694 43488 5702 43552
rect 5382 42464 5702 43488
rect 5382 42400 5390 42464
rect 5454 42400 5470 42464
rect 5534 42400 5550 42464
rect 5614 42400 5630 42464
rect 5694 42400 5702 42464
rect 5382 41376 5702 42400
rect 5382 41312 5390 41376
rect 5454 41312 5470 41376
rect 5534 41312 5550 41376
rect 5614 41312 5630 41376
rect 5694 41312 5702 41376
rect 5382 40288 5702 41312
rect 5382 40224 5390 40288
rect 5454 40224 5470 40288
rect 5534 40224 5550 40288
rect 5614 40224 5630 40288
rect 5694 40224 5702 40288
rect 5382 39200 5702 40224
rect 5382 39136 5390 39200
rect 5454 39136 5470 39200
rect 5534 39136 5550 39200
rect 5614 39136 5630 39200
rect 5694 39136 5702 39200
rect 5382 38112 5702 39136
rect 5382 38048 5390 38112
rect 5454 38048 5470 38112
rect 5534 38048 5550 38112
rect 5614 38048 5630 38112
rect 5694 38048 5702 38112
rect 5382 37024 5702 38048
rect 5382 36960 5390 37024
rect 5454 36960 5470 37024
rect 5534 36960 5550 37024
rect 5614 36960 5630 37024
rect 5694 36960 5702 37024
rect 5382 35936 5702 36960
rect 5382 35872 5390 35936
rect 5454 35872 5470 35936
rect 5534 35872 5550 35936
rect 5614 35872 5630 35936
rect 5694 35872 5702 35936
rect 5382 34848 5702 35872
rect 5382 34784 5390 34848
rect 5454 34784 5470 34848
rect 5534 34784 5550 34848
rect 5614 34784 5630 34848
rect 5694 34784 5702 34848
rect 5382 33760 5702 34784
rect 5382 33696 5390 33760
rect 5454 33696 5470 33760
rect 5534 33696 5550 33760
rect 5614 33696 5630 33760
rect 5694 33696 5702 33760
rect 5382 32672 5702 33696
rect 5382 32608 5390 32672
rect 5454 32608 5470 32672
rect 5534 32608 5550 32672
rect 5614 32608 5630 32672
rect 5694 32608 5702 32672
rect 5382 31584 5702 32608
rect 5382 31520 5390 31584
rect 5454 31520 5470 31584
rect 5534 31520 5550 31584
rect 5614 31520 5630 31584
rect 5694 31520 5702 31584
rect 5382 30496 5702 31520
rect 5382 30432 5390 30496
rect 5454 30432 5470 30496
rect 5534 30432 5550 30496
rect 5614 30432 5630 30496
rect 5694 30432 5702 30496
rect 4659 30428 4725 30429
rect 4659 30364 4660 30428
rect 4724 30364 4725 30428
rect 4659 30363 4725 30364
rect 3163 29888 3171 29952
rect 3235 29888 3251 29952
rect 3315 29888 3331 29952
rect 3395 29888 3411 29952
rect 3475 29888 3483 29952
rect 3163 28864 3483 29888
rect 3163 28800 3171 28864
rect 3235 28800 3251 28864
rect 3315 28800 3331 28864
rect 3395 28800 3411 28864
rect 3475 28800 3483 28864
rect 3163 27776 3483 28800
rect 3163 27712 3171 27776
rect 3235 27712 3251 27776
rect 3315 27712 3331 27776
rect 3395 27712 3411 27776
rect 3475 27712 3483 27776
rect 3163 26688 3483 27712
rect 4291 27708 4357 27709
rect 4291 27644 4292 27708
rect 4356 27644 4357 27708
rect 4291 27643 4357 27644
rect 3163 26624 3171 26688
rect 3235 26624 3251 26688
rect 3315 26624 3331 26688
rect 3395 26624 3411 26688
rect 3475 26624 3483 26688
rect 1899 26620 1965 26621
rect 1899 26556 1900 26620
rect 1964 26556 1965 26620
rect 1899 26555 1965 26556
rect 1902 11661 1962 26555
rect 3163 25600 3483 26624
rect 3163 25536 3171 25600
rect 3235 25536 3251 25600
rect 3315 25536 3331 25600
rect 3395 25536 3411 25600
rect 3475 25536 3483 25600
rect 3163 24512 3483 25536
rect 3163 24448 3171 24512
rect 3235 24448 3251 24512
rect 3315 24448 3331 24512
rect 3395 24448 3411 24512
rect 3475 24448 3483 24512
rect 3163 23424 3483 24448
rect 3923 23492 3989 23493
rect 3923 23428 3924 23492
rect 3988 23428 3989 23492
rect 3923 23427 3989 23428
rect 3163 23360 3171 23424
rect 3235 23360 3251 23424
rect 3315 23360 3331 23424
rect 3395 23360 3411 23424
rect 3475 23360 3483 23424
rect 3163 22336 3483 23360
rect 3163 22272 3171 22336
rect 3235 22272 3251 22336
rect 3315 22272 3331 22336
rect 3395 22272 3411 22336
rect 3475 22272 3483 22336
rect 3163 21248 3483 22272
rect 3163 21184 3171 21248
rect 3235 21184 3251 21248
rect 3315 21184 3331 21248
rect 3395 21184 3411 21248
rect 3475 21184 3483 21248
rect 3163 20160 3483 21184
rect 3163 20096 3171 20160
rect 3235 20096 3251 20160
rect 3315 20096 3331 20160
rect 3395 20096 3411 20160
rect 3475 20096 3483 20160
rect 2083 19412 2149 19413
rect 2083 19348 2084 19412
rect 2148 19348 2149 19412
rect 2083 19347 2149 19348
rect 2086 13837 2146 19347
rect 3163 19072 3483 20096
rect 3163 19008 3171 19072
rect 3235 19008 3251 19072
rect 3315 19008 3331 19072
rect 3395 19008 3411 19072
rect 3475 19008 3483 19072
rect 3163 17984 3483 19008
rect 3163 17920 3171 17984
rect 3235 17920 3251 17984
rect 3315 17920 3331 17984
rect 3395 17920 3411 17984
rect 3475 17920 3483 17984
rect 3163 16896 3483 17920
rect 3926 17237 3986 23427
rect 3923 17236 3989 17237
rect 3923 17172 3924 17236
rect 3988 17172 3989 17236
rect 3923 17171 3989 17172
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3003 16692 3069 16693
rect 3003 16628 3004 16692
rect 3068 16628 3069 16692
rect 3003 16627 3069 16628
rect 2083 13836 2149 13837
rect 2083 13772 2084 13836
rect 2148 13772 2149 13836
rect 2083 13771 2149 13772
rect 1899 11660 1965 11661
rect 1899 11596 1900 11660
rect 1964 11596 1965 11660
rect 1899 11595 1965 11596
rect 3006 9757 3066 16627
rect 3163 15808 3483 16832
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 14720 3483 15744
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3163 13632 3483 14656
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11456 3483 12480
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 4294 10981 4354 27643
rect 4291 10980 4357 10981
rect 4291 10916 4292 10980
rect 4356 10916 4357 10980
rect 4291 10915 4357 10916
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3003 9756 3069 9757
rect 3003 9692 3004 9756
rect 3068 9692 3069 9756
rect 3003 9691 3069 9692
rect 3163 9280 3483 10304
rect 4662 9621 4722 30363
rect 5382 29408 5702 30432
rect 5382 29344 5390 29408
rect 5454 29344 5470 29408
rect 5534 29344 5550 29408
rect 5614 29344 5630 29408
rect 5694 29344 5702 29408
rect 5382 28320 5702 29344
rect 5382 28256 5390 28320
rect 5454 28256 5470 28320
rect 5534 28256 5550 28320
rect 5614 28256 5630 28320
rect 5694 28256 5702 28320
rect 5382 27232 5702 28256
rect 5382 27168 5390 27232
rect 5454 27168 5470 27232
rect 5534 27168 5550 27232
rect 5614 27168 5630 27232
rect 5694 27168 5702 27232
rect 5382 26144 5702 27168
rect 7602 47360 7922 47376
rect 7602 47296 7610 47360
rect 7674 47296 7690 47360
rect 7754 47296 7770 47360
rect 7834 47296 7850 47360
rect 7914 47296 7922 47360
rect 7602 46272 7922 47296
rect 7602 46208 7610 46272
rect 7674 46208 7690 46272
rect 7754 46208 7770 46272
rect 7834 46208 7850 46272
rect 7914 46208 7922 46272
rect 7602 45184 7922 46208
rect 7602 45120 7610 45184
rect 7674 45120 7690 45184
rect 7754 45120 7770 45184
rect 7834 45120 7850 45184
rect 7914 45120 7922 45184
rect 7602 44096 7922 45120
rect 7602 44032 7610 44096
rect 7674 44032 7690 44096
rect 7754 44032 7770 44096
rect 7834 44032 7850 44096
rect 7914 44032 7922 44096
rect 7602 43008 7922 44032
rect 7602 42944 7610 43008
rect 7674 42944 7690 43008
rect 7754 42944 7770 43008
rect 7834 42944 7850 43008
rect 7914 42944 7922 43008
rect 7602 41920 7922 42944
rect 7602 41856 7610 41920
rect 7674 41856 7690 41920
rect 7754 41856 7770 41920
rect 7834 41856 7850 41920
rect 7914 41856 7922 41920
rect 7602 40832 7922 41856
rect 7602 40768 7610 40832
rect 7674 40768 7690 40832
rect 7754 40768 7770 40832
rect 7834 40768 7850 40832
rect 7914 40768 7922 40832
rect 7602 39744 7922 40768
rect 7602 39680 7610 39744
rect 7674 39680 7690 39744
rect 7754 39680 7770 39744
rect 7834 39680 7850 39744
rect 7914 39680 7922 39744
rect 7602 38656 7922 39680
rect 7602 38592 7610 38656
rect 7674 38592 7690 38656
rect 7754 38592 7770 38656
rect 7834 38592 7850 38656
rect 7914 38592 7922 38656
rect 7602 37568 7922 38592
rect 7602 37504 7610 37568
rect 7674 37504 7690 37568
rect 7754 37504 7770 37568
rect 7834 37504 7850 37568
rect 7914 37504 7922 37568
rect 7602 36480 7922 37504
rect 7602 36416 7610 36480
rect 7674 36416 7690 36480
rect 7754 36416 7770 36480
rect 7834 36416 7850 36480
rect 7914 36416 7922 36480
rect 7602 35392 7922 36416
rect 7602 35328 7610 35392
rect 7674 35328 7690 35392
rect 7754 35328 7770 35392
rect 7834 35328 7850 35392
rect 7914 35328 7922 35392
rect 7602 34304 7922 35328
rect 7602 34240 7610 34304
rect 7674 34240 7690 34304
rect 7754 34240 7770 34304
rect 7834 34240 7850 34304
rect 7914 34240 7922 34304
rect 7602 33216 7922 34240
rect 7602 33152 7610 33216
rect 7674 33152 7690 33216
rect 7754 33152 7770 33216
rect 7834 33152 7850 33216
rect 7914 33152 7922 33216
rect 7602 32128 7922 33152
rect 7602 32064 7610 32128
rect 7674 32064 7690 32128
rect 7754 32064 7770 32128
rect 7834 32064 7850 32128
rect 7914 32064 7922 32128
rect 7602 31040 7922 32064
rect 7602 30976 7610 31040
rect 7674 30976 7690 31040
rect 7754 30976 7770 31040
rect 7834 30976 7850 31040
rect 7914 30976 7922 31040
rect 7602 29952 7922 30976
rect 7602 29888 7610 29952
rect 7674 29888 7690 29952
rect 7754 29888 7770 29952
rect 7834 29888 7850 29952
rect 7914 29888 7922 29952
rect 7602 28864 7922 29888
rect 9821 46816 10141 47376
rect 9821 46752 9829 46816
rect 9893 46752 9909 46816
rect 9973 46752 9989 46816
rect 10053 46752 10069 46816
rect 10133 46752 10141 46816
rect 9821 45728 10141 46752
rect 9821 45664 9829 45728
rect 9893 45664 9909 45728
rect 9973 45664 9989 45728
rect 10053 45664 10069 45728
rect 10133 45664 10141 45728
rect 9821 44640 10141 45664
rect 9821 44576 9829 44640
rect 9893 44576 9909 44640
rect 9973 44576 9989 44640
rect 10053 44576 10069 44640
rect 10133 44576 10141 44640
rect 9821 43552 10141 44576
rect 9821 43488 9829 43552
rect 9893 43488 9909 43552
rect 9973 43488 9989 43552
rect 10053 43488 10069 43552
rect 10133 43488 10141 43552
rect 9821 42464 10141 43488
rect 9821 42400 9829 42464
rect 9893 42400 9909 42464
rect 9973 42400 9989 42464
rect 10053 42400 10069 42464
rect 10133 42400 10141 42464
rect 9821 41376 10141 42400
rect 9821 41312 9829 41376
rect 9893 41312 9909 41376
rect 9973 41312 9989 41376
rect 10053 41312 10069 41376
rect 10133 41312 10141 41376
rect 9821 40288 10141 41312
rect 9821 40224 9829 40288
rect 9893 40224 9909 40288
rect 9973 40224 9989 40288
rect 10053 40224 10069 40288
rect 10133 40224 10141 40288
rect 9821 39200 10141 40224
rect 9821 39136 9829 39200
rect 9893 39136 9909 39200
rect 9973 39136 9989 39200
rect 10053 39136 10069 39200
rect 10133 39136 10141 39200
rect 9821 38112 10141 39136
rect 9821 38048 9829 38112
rect 9893 38048 9909 38112
rect 9973 38048 9989 38112
rect 10053 38048 10069 38112
rect 10133 38048 10141 38112
rect 9821 37024 10141 38048
rect 9821 36960 9829 37024
rect 9893 36960 9909 37024
rect 9973 36960 9989 37024
rect 10053 36960 10069 37024
rect 10133 36960 10141 37024
rect 9821 35936 10141 36960
rect 9821 35872 9829 35936
rect 9893 35872 9909 35936
rect 9973 35872 9989 35936
rect 10053 35872 10069 35936
rect 10133 35872 10141 35936
rect 9821 34848 10141 35872
rect 9821 34784 9829 34848
rect 9893 34784 9909 34848
rect 9973 34784 9989 34848
rect 10053 34784 10069 34848
rect 10133 34784 10141 34848
rect 9821 33760 10141 34784
rect 9821 33696 9829 33760
rect 9893 33696 9909 33760
rect 9973 33696 9989 33760
rect 10053 33696 10069 33760
rect 10133 33696 10141 33760
rect 9821 32672 10141 33696
rect 9821 32608 9829 32672
rect 9893 32608 9909 32672
rect 9973 32608 9989 32672
rect 10053 32608 10069 32672
rect 10133 32608 10141 32672
rect 9821 31584 10141 32608
rect 9821 31520 9829 31584
rect 9893 31520 9909 31584
rect 9973 31520 9989 31584
rect 10053 31520 10069 31584
rect 10133 31520 10141 31584
rect 9821 30496 10141 31520
rect 9821 30432 9829 30496
rect 9893 30432 9909 30496
rect 9973 30432 9989 30496
rect 10053 30432 10069 30496
rect 10133 30432 10141 30496
rect 9821 29408 10141 30432
rect 9821 29344 9829 29408
rect 9893 29344 9909 29408
rect 9973 29344 9989 29408
rect 10053 29344 10069 29408
rect 10133 29344 10141 29408
rect 8155 29068 8221 29069
rect 8155 29004 8156 29068
rect 8220 29004 8221 29068
rect 8155 29003 8221 29004
rect 7602 28800 7610 28864
rect 7674 28800 7690 28864
rect 7754 28800 7770 28864
rect 7834 28800 7850 28864
rect 7914 28800 7922 28864
rect 7602 27776 7922 28800
rect 7602 27712 7610 27776
rect 7674 27712 7690 27776
rect 7754 27712 7770 27776
rect 7834 27712 7850 27776
rect 7914 27712 7922 27776
rect 7419 27164 7485 27165
rect 7419 27100 7420 27164
rect 7484 27100 7485 27164
rect 7419 27099 7485 27100
rect 6683 26348 6749 26349
rect 6683 26284 6684 26348
rect 6748 26284 6749 26348
rect 6683 26283 6749 26284
rect 5382 26080 5390 26144
rect 5454 26080 5470 26144
rect 5534 26080 5550 26144
rect 5614 26080 5630 26144
rect 5694 26080 5702 26144
rect 4843 25260 4909 25261
rect 4843 25196 4844 25260
rect 4908 25196 4909 25260
rect 4843 25195 4909 25196
rect 4659 9620 4725 9621
rect 4659 9556 4660 9620
rect 4724 9556 4725 9620
rect 4659 9555 4725 9556
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 7104 3483 8128
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 4846 5541 4906 25195
rect 5382 25056 5702 26080
rect 5382 24992 5390 25056
rect 5454 24992 5470 25056
rect 5534 24992 5550 25056
rect 5614 24992 5630 25056
rect 5694 24992 5702 25056
rect 5382 23968 5702 24992
rect 5382 23904 5390 23968
rect 5454 23904 5470 23968
rect 5534 23904 5550 23968
rect 5614 23904 5630 23968
rect 5694 23904 5702 23968
rect 5382 22880 5702 23904
rect 5382 22816 5390 22880
rect 5454 22816 5470 22880
rect 5534 22816 5550 22880
rect 5614 22816 5630 22880
rect 5694 22816 5702 22880
rect 5382 21792 5702 22816
rect 5382 21728 5390 21792
rect 5454 21728 5470 21792
rect 5534 21728 5550 21792
rect 5614 21728 5630 21792
rect 5694 21728 5702 21792
rect 5382 20704 5702 21728
rect 5382 20640 5390 20704
rect 5454 20640 5470 20704
rect 5534 20640 5550 20704
rect 5614 20640 5630 20704
rect 5694 20640 5702 20704
rect 5382 19616 5702 20640
rect 5382 19552 5390 19616
rect 5454 19552 5470 19616
rect 5534 19552 5550 19616
rect 5614 19552 5630 19616
rect 5694 19552 5702 19616
rect 5382 18528 5702 19552
rect 5382 18464 5390 18528
rect 5454 18464 5470 18528
rect 5534 18464 5550 18528
rect 5614 18464 5630 18528
rect 5694 18464 5702 18528
rect 5382 17440 5702 18464
rect 5382 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5702 17440
rect 5382 16352 5702 17376
rect 5382 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5702 16352
rect 5382 15264 5702 16288
rect 5382 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5702 15264
rect 5382 14176 5702 15200
rect 5382 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5702 14176
rect 5382 13088 5702 14112
rect 5382 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5702 13088
rect 5382 12000 5702 13024
rect 5382 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5702 12000
rect 5382 10912 5702 11936
rect 5382 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5702 10912
rect 5382 9824 5702 10848
rect 5382 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5702 9824
rect 5382 8736 5702 9760
rect 5382 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5702 8736
rect 5382 7648 5702 8672
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 6686 6629 6746 26283
rect 7422 24173 7482 27099
rect 7602 26688 7922 27712
rect 7602 26624 7610 26688
rect 7674 26624 7690 26688
rect 7754 26624 7770 26688
rect 7834 26624 7850 26688
rect 7914 26624 7922 26688
rect 7602 25600 7922 26624
rect 7602 25536 7610 25600
rect 7674 25536 7690 25600
rect 7754 25536 7770 25600
rect 7834 25536 7850 25600
rect 7914 25536 7922 25600
rect 7602 24512 7922 25536
rect 7602 24448 7610 24512
rect 7674 24448 7690 24512
rect 7754 24448 7770 24512
rect 7834 24448 7850 24512
rect 7914 24448 7922 24512
rect 7419 24172 7485 24173
rect 7419 24108 7420 24172
rect 7484 24108 7485 24172
rect 7419 24107 7485 24108
rect 7602 23424 7922 24448
rect 7602 23360 7610 23424
rect 7674 23360 7690 23424
rect 7754 23360 7770 23424
rect 7834 23360 7850 23424
rect 7914 23360 7922 23424
rect 7602 22336 7922 23360
rect 7602 22272 7610 22336
rect 7674 22272 7690 22336
rect 7754 22272 7770 22336
rect 7834 22272 7850 22336
rect 7914 22272 7922 22336
rect 7602 21248 7922 22272
rect 7602 21184 7610 21248
rect 7674 21184 7690 21248
rect 7754 21184 7770 21248
rect 7834 21184 7850 21248
rect 7914 21184 7922 21248
rect 7602 20160 7922 21184
rect 8158 20773 8218 29003
rect 9821 28320 10141 29344
rect 9821 28256 9829 28320
rect 9893 28256 9909 28320
rect 9973 28256 9989 28320
rect 10053 28256 10069 28320
rect 10133 28256 10141 28320
rect 9821 27232 10141 28256
rect 9821 27168 9829 27232
rect 9893 27168 9909 27232
rect 9973 27168 9989 27232
rect 10053 27168 10069 27232
rect 10133 27168 10141 27232
rect 9821 26144 10141 27168
rect 9821 26080 9829 26144
rect 9893 26080 9909 26144
rect 9973 26080 9989 26144
rect 10053 26080 10069 26144
rect 10133 26080 10141 26144
rect 9821 25056 10141 26080
rect 9821 24992 9829 25056
rect 9893 24992 9909 25056
rect 9973 24992 9989 25056
rect 10053 24992 10069 25056
rect 10133 24992 10141 25056
rect 9821 23968 10141 24992
rect 9821 23904 9829 23968
rect 9893 23904 9909 23968
rect 9973 23904 9989 23968
rect 10053 23904 10069 23968
rect 10133 23904 10141 23968
rect 9821 22880 10141 23904
rect 9821 22816 9829 22880
rect 9893 22816 9909 22880
rect 9973 22816 9989 22880
rect 10053 22816 10069 22880
rect 10133 22816 10141 22880
rect 9821 21792 10141 22816
rect 9821 21728 9829 21792
rect 9893 21728 9909 21792
rect 9973 21728 9989 21792
rect 10053 21728 10069 21792
rect 10133 21728 10141 21792
rect 8155 20772 8221 20773
rect 8155 20708 8156 20772
rect 8220 20708 8221 20772
rect 8155 20707 8221 20708
rect 7602 20096 7610 20160
rect 7674 20096 7690 20160
rect 7754 20096 7770 20160
rect 7834 20096 7850 20160
rect 7914 20096 7922 20160
rect 7602 19072 7922 20096
rect 7602 19008 7610 19072
rect 7674 19008 7690 19072
rect 7754 19008 7770 19072
rect 7834 19008 7850 19072
rect 7914 19008 7922 19072
rect 7602 17984 7922 19008
rect 7602 17920 7610 17984
rect 7674 17920 7690 17984
rect 7754 17920 7770 17984
rect 7834 17920 7850 17984
rect 7914 17920 7922 17984
rect 7602 16896 7922 17920
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 7602 15808 7922 16832
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 14720 7922 15744
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7602 11456 7922 12480
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7602 9280 7922 10304
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 7602 7104 7922 8128
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 6683 6628 6749 6629
rect 6683 6564 6684 6628
rect 6748 6564 6749 6628
rect 6683 6563 6749 6564
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 4843 5540 4909 5541
rect 4843 5476 4844 5540
rect 4908 5476 4909 5540
rect 4843 5475 4909 5476
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 20704 10141 21728
rect 9821 20640 9829 20704
rect 9893 20640 9909 20704
rect 9973 20640 9989 20704
rect 10053 20640 10069 20704
rect 10133 20640 10141 20704
rect 9821 19616 10141 20640
rect 9821 19552 9829 19616
rect 9893 19552 9909 19616
rect 9973 19552 9989 19616
rect 10053 19552 10069 19616
rect 10133 19552 10141 19616
rect 9821 18528 10141 19552
rect 9821 18464 9829 18528
rect 9893 18464 9909 18528
rect 9973 18464 9989 18528
rect 10053 18464 10069 18528
rect 10133 18464 10141 18528
rect 9821 17440 10141 18464
rect 9821 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10141 17440
rect 9821 16352 10141 17376
rect 9821 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10141 16352
rect 9821 15264 10141 16288
rect 9821 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10141 15264
rect 9821 14176 10141 15200
rect 9821 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10141 14176
rect 9821 13088 10141 14112
rect 9821 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10141 13088
rect 9821 12000 10141 13024
rect 9821 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10141 12000
rect 9821 10912 10141 11936
rect 9821 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10141 10912
rect 9821 9824 10141 10848
rect 9821 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10141 9824
rect 9821 8736 10141 9760
rect 9821 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10141 8736
rect 9821 7648 10141 8672
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 47360 12361 47376
rect 12041 47296 12049 47360
rect 12113 47296 12129 47360
rect 12193 47296 12209 47360
rect 12273 47296 12289 47360
rect 12353 47296 12361 47360
rect 12041 46272 12361 47296
rect 12041 46208 12049 46272
rect 12113 46208 12129 46272
rect 12193 46208 12209 46272
rect 12273 46208 12289 46272
rect 12353 46208 12361 46272
rect 12041 45184 12361 46208
rect 12041 45120 12049 45184
rect 12113 45120 12129 45184
rect 12193 45120 12209 45184
rect 12273 45120 12289 45184
rect 12353 45120 12361 45184
rect 12041 44096 12361 45120
rect 12041 44032 12049 44096
rect 12113 44032 12129 44096
rect 12193 44032 12209 44096
rect 12273 44032 12289 44096
rect 12353 44032 12361 44096
rect 12041 43008 12361 44032
rect 12041 42944 12049 43008
rect 12113 42944 12129 43008
rect 12193 42944 12209 43008
rect 12273 42944 12289 43008
rect 12353 42944 12361 43008
rect 12041 41920 12361 42944
rect 12041 41856 12049 41920
rect 12113 41856 12129 41920
rect 12193 41856 12209 41920
rect 12273 41856 12289 41920
rect 12353 41856 12361 41920
rect 12041 40832 12361 41856
rect 12041 40768 12049 40832
rect 12113 40768 12129 40832
rect 12193 40768 12209 40832
rect 12273 40768 12289 40832
rect 12353 40768 12361 40832
rect 12041 39744 12361 40768
rect 12041 39680 12049 39744
rect 12113 39680 12129 39744
rect 12193 39680 12209 39744
rect 12273 39680 12289 39744
rect 12353 39680 12361 39744
rect 12041 38656 12361 39680
rect 12041 38592 12049 38656
rect 12113 38592 12129 38656
rect 12193 38592 12209 38656
rect 12273 38592 12289 38656
rect 12353 38592 12361 38656
rect 12041 37568 12361 38592
rect 12041 37504 12049 37568
rect 12113 37504 12129 37568
rect 12193 37504 12209 37568
rect 12273 37504 12289 37568
rect 12353 37504 12361 37568
rect 12041 36480 12361 37504
rect 12041 36416 12049 36480
rect 12113 36416 12129 36480
rect 12193 36416 12209 36480
rect 12273 36416 12289 36480
rect 12353 36416 12361 36480
rect 12041 35392 12361 36416
rect 12041 35328 12049 35392
rect 12113 35328 12129 35392
rect 12193 35328 12209 35392
rect 12273 35328 12289 35392
rect 12353 35328 12361 35392
rect 12041 34304 12361 35328
rect 12041 34240 12049 34304
rect 12113 34240 12129 34304
rect 12193 34240 12209 34304
rect 12273 34240 12289 34304
rect 12353 34240 12361 34304
rect 12041 33216 12361 34240
rect 12041 33152 12049 33216
rect 12113 33152 12129 33216
rect 12193 33152 12209 33216
rect 12273 33152 12289 33216
rect 12353 33152 12361 33216
rect 12041 32128 12361 33152
rect 12041 32064 12049 32128
rect 12113 32064 12129 32128
rect 12193 32064 12209 32128
rect 12273 32064 12289 32128
rect 12353 32064 12361 32128
rect 12041 31040 12361 32064
rect 12041 30976 12049 31040
rect 12113 30976 12129 31040
rect 12193 30976 12209 31040
rect 12273 30976 12289 31040
rect 12353 30976 12361 31040
rect 12041 29952 12361 30976
rect 12041 29888 12049 29952
rect 12113 29888 12129 29952
rect 12193 29888 12209 29952
rect 12273 29888 12289 29952
rect 12353 29888 12361 29952
rect 12041 28864 12361 29888
rect 12041 28800 12049 28864
rect 12113 28800 12129 28864
rect 12193 28800 12209 28864
rect 12273 28800 12289 28864
rect 12353 28800 12361 28864
rect 12041 27776 12361 28800
rect 12041 27712 12049 27776
rect 12113 27712 12129 27776
rect 12193 27712 12209 27776
rect 12273 27712 12289 27776
rect 12353 27712 12361 27776
rect 12041 26688 12361 27712
rect 12041 26624 12049 26688
rect 12113 26624 12129 26688
rect 12193 26624 12209 26688
rect 12273 26624 12289 26688
rect 12353 26624 12361 26688
rect 12041 25600 12361 26624
rect 12041 25536 12049 25600
rect 12113 25536 12129 25600
rect 12193 25536 12209 25600
rect 12273 25536 12289 25600
rect 12353 25536 12361 25600
rect 12041 24512 12361 25536
rect 12041 24448 12049 24512
rect 12113 24448 12129 24512
rect 12193 24448 12209 24512
rect 12273 24448 12289 24512
rect 12353 24448 12361 24512
rect 12041 23424 12361 24448
rect 12041 23360 12049 23424
rect 12113 23360 12129 23424
rect 12193 23360 12209 23424
rect 12273 23360 12289 23424
rect 12353 23360 12361 23424
rect 12041 22336 12361 23360
rect 12041 22272 12049 22336
rect 12113 22272 12129 22336
rect 12193 22272 12209 22336
rect 12273 22272 12289 22336
rect 12353 22272 12361 22336
rect 12041 21248 12361 22272
rect 12041 21184 12049 21248
rect 12113 21184 12129 21248
rect 12193 21184 12209 21248
rect 12273 21184 12289 21248
rect 12353 21184 12361 21248
rect 12041 20160 12361 21184
rect 12041 20096 12049 20160
rect 12113 20096 12129 20160
rect 12193 20096 12209 20160
rect 12273 20096 12289 20160
rect 12353 20096 12361 20160
rect 12041 19072 12361 20096
rect 12041 19008 12049 19072
rect 12113 19008 12129 19072
rect 12193 19008 12209 19072
rect 12273 19008 12289 19072
rect 12353 19008 12361 19072
rect 12041 17984 12361 19008
rect 12041 17920 12049 17984
rect 12113 17920 12129 17984
rect 12193 17920 12209 17984
rect 12273 17920 12289 17984
rect 12353 17920 12361 17984
rect 12041 16896 12361 17920
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 12041 14720 12361 15744
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 12041 13632 12361 14656
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 12041 11456 12361 12480
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 12041 9280 12361 10304
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 7104 12361 8128
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 46816 14580 47376
rect 14260 46752 14268 46816
rect 14332 46752 14348 46816
rect 14412 46752 14428 46816
rect 14492 46752 14508 46816
rect 14572 46752 14580 46816
rect 14260 45728 14580 46752
rect 14260 45664 14268 45728
rect 14332 45664 14348 45728
rect 14412 45664 14428 45728
rect 14492 45664 14508 45728
rect 14572 45664 14580 45728
rect 14260 44640 14580 45664
rect 14260 44576 14268 44640
rect 14332 44576 14348 44640
rect 14412 44576 14428 44640
rect 14492 44576 14508 44640
rect 14572 44576 14580 44640
rect 14260 43552 14580 44576
rect 14260 43488 14268 43552
rect 14332 43488 14348 43552
rect 14412 43488 14428 43552
rect 14492 43488 14508 43552
rect 14572 43488 14580 43552
rect 14260 42464 14580 43488
rect 14260 42400 14268 42464
rect 14332 42400 14348 42464
rect 14412 42400 14428 42464
rect 14492 42400 14508 42464
rect 14572 42400 14580 42464
rect 14260 41376 14580 42400
rect 14260 41312 14268 41376
rect 14332 41312 14348 41376
rect 14412 41312 14428 41376
rect 14492 41312 14508 41376
rect 14572 41312 14580 41376
rect 14260 40288 14580 41312
rect 14260 40224 14268 40288
rect 14332 40224 14348 40288
rect 14412 40224 14428 40288
rect 14492 40224 14508 40288
rect 14572 40224 14580 40288
rect 14260 39200 14580 40224
rect 14260 39136 14268 39200
rect 14332 39136 14348 39200
rect 14412 39136 14428 39200
rect 14492 39136 14508 39200
rect 14572 39136 14580 39200
rect 14260 38112 14580 39136
rect 14260 38048 14268 38112
rect 14332 38048 14348 38112
rect 14412 38048 14428 38112
rect 14492 38048 14508 38112
rect 14572 38048 14580 38112
rect 14260 37024 14580 38048
rect 14260 36960 14268 37024
rect 14332 36960 14348 37024
rect 14412 36960 14428 37024
rect 14492 36960 14508 37024
rect 14572 36960 14580 37024
rect 14260 35936 14580 36960
rect 14260 35872 14268 35936
rect 14332 35872 14348 35936
rect 14412 35872 14428 35936
rect 14492 35872 14508 35936
rect 14572 35872 14580 35936
rect 14260 34848 14580 35872
rect 14260 34784 14268 34848
rect 14332 34784 14348 34848
rect 14412 34784 14428 34848
rect 14492 34784 14508 34848
rect 14572 34784 14580 34848
rect 14260 33760 14580 34784
rect 14260 33696 14268 33760
rect 14332 33696 14348 33760
rect 14412 33696 14428 33760
rect 14492 33696 14508 33760
rect 14572 33696 14580 33760
rect 14260 32672 14580 33696
rect 14260 32608 14268 32672
rect 14332 32608 14348 32672
rect 14412 32608 14428 32672
rect 14492 32608 14508 32672
rect 14572 32608 14580 32672
rect 14260 31584 14580 32608
rect 14260 31520 14268 31584
rect 14332 31520 14348 31584
rect 14412 31520 14428 31584
rect 14492 31520 14508 31584
rect 14572 31520 14580 31584
rect 14260 30496 14580 31520
rect 14260 30432 14268 30496
rect 14332 30432 14348 30496
rect 14412 30432 14428 30496
rect 14492 30432 14508 30496
rect 14572 30432 14580 30496
rect 14260 29408 14580 30432
rect 14260 29344 14268 29408
rect 14332 29344 14348 29408
rect 14412 29344 14428 29408
rect 14492 29344 14508 29408
rect 14572 29344 14580 29408
rect 14260 28320 14580 29344
rect 14260 28256 14268 28320
rect 14332 28256 14348 28320
rect 14412 28256 14428 28320
rect 14492 28256 14508 28320
rect 14572 28256 14580 28320
rect 14260 27232 14580 28256
rect 14260 27168 14268 27232
rect 14332 27168 14348 27232
rect 14412 27168 14428 27232
rect 14492 27168 14508 27232
rect 14572 27168 14580 27232
rect 14260 26144 14580 27168
rect 14260 26080 14268 26144
rect 14332 26080 14348 26144
rect 14412 26080 14428 26144
rect 14492 26080 14508 26144
rect 14572 26080 14580 26144
rect 14260 25056 14580 26080
rect 14260 24992 14268 25056
rect 14332 24992 14348 25056
rect 14412 24992 14428 25056
rect 14492 24992 14508 25056
rect 14572 24992 14580 25056
rect 14260 23968 14580 24992
rect 14260 23904 14268 23968
rect 14332 23904 14348 23968
rect 14412 23904 14428 23968
rect 14492 23904 14508 23968
rect 14572 23904 14580 23968
rect 14260 22880 14580 23904
rect 14260 22816 14268 22880
rect 14332 22816 14348 22880
rect 14412 22816 14428 22880
rect 14492 22816 14508 22880
rect 14572 22816 14580 22880
rect 14260 21792 14580 22816
rect 14260 21728 14268 21792
rect 14332 21728 14348 21792
rect 14412 21728 14428 21792
rect 14492 21728 14508 21792
rect 14572 21728 14580 21792
rect 14260 20704 14580 21728
rect 14260 20640 14268 20704
rect 14332 20640 14348 20704
rect 14412 20640 14428 20704
rect 14492 20640 14508 20704
rect 14572 20640 14580 20704
rect 14260 19616 14580 20640
rect 14260 19552 14268 19616
rect 14332 19552 14348 19616
rect 14412 19552 14428 19616
rect 14492 19552 14508 19616
rect 14572 19552 14580 19616
rect 14260 18528 14580 19552
rect 14260 18464 14268 18528
rect 14332 18464 14348 18528
rect 14412 18464 14428 18528
rect 14492 18464 14508 18528
rect 14572 18464 14580 18528
rect 14260 17440 14580 18464
rect 14260 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14580 17440
rect 14260 16352 14580 17376
rect 14260 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14580 16352
rect 14260 15264 14580 16288
rect 14260 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14580 15264
rect 14260 14176 14580 15200
rect 14260 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14580 14176
rect 14260 13088 14580 14112
rect 14260 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14580 13088
rect 14260 12000 14580 13024
rect 14260 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14580 12000
rect 14260 10912 14580 11936
rect 14260 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14580 10912
rect 14260 9824 14580 10848
rect 14260 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14580 9824
rect 14260 8736 14580 9760
rect 14260 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14580 8736
rect 14260 7648 14580 8672
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 47360 16800 47376
rect 16480 47296 16488 47360
rect 16552 47296 16568 47360
rect 16632 47296 16648 47360
rect 16712 47296 16728 47360
rect 16792 47296 16800 47360
rect 16480 46272 16800 47296
rect 16480 46208 16488 46272
rect 16552 46208 16568 46272
rect 16632 46208 16648 46272
rect 16712 46208 16728 46272
rect 16792 46208 16800 46272
rect 16480 45184 16800 46208
rect 16480 45120 16488 45184
rect 16552 45120 16568 45184
rect 16632 45120 16648 45184
rect 16712 45120 16728 45184
rect 16792 45120 16800 45184
rect 16480 44096 16800 45120
rect 16480 44032 16488 44096
rect 16552 44032 16568 44096
rect 16632 44032 16648 44096
rect 16712 44032 16728 44096
rect 16792 44032 16800 44096
rect 16480 43008 16800 44032
rect 16480 42944 16488 43008
rect 16552 42944 16568 43008
rect 16632 42944 16648 43008
rect 16712 42944 16728 43008
rect 16792 42944 16800 43008
rect 16480 41920 16800 42944
rect 16480 41856 16488 41920
rect 16552 41856 16568 41920
rect 16632 41856 16648 41920
rect 16712 41856 16728 41920
rect 16792 41856 16800 41920
rect 16480 40832 16800 41856
rect 16480 40768 16488 40832
rect 16552 40768 16568 40832
rect 16632 40768 16648 40832
rect 16712 40768 16728 40832
rect 16792 40768 16800 40832
rect 16480 39744 16800 40768
rect 16480 39680 16488 39744
rect 16552 39680 16568 39744
rect 16632 39680 16648 39744
rect 16712 39680 16728 39744
rect 16792 39680 16800 39744
rect 16480 38656 16800 39680
rect 16480 38592 16488 38656
rect 16552 38592 16568 38656
rect 16632 38592 16648 38656
rect 16712 38592 16728 38656
rect 16792 38592 16800 38656
rect 16480 37568 16800 38592
rect 16480 37504 16488 37568
rect 16552 37504 16568 37568
rect 16632 37504 16648 37568
rect 16712 37504 16728 37568
rect 16792 37504 16800 37568
rect 16480 36480 16800 37504
rect 16480 36416 16488 36480
rect 16552 36416 16568 36480
rect 16632 36416 16648 36480
rect 16712 36416 16728 36480
rect 16792 36416 16800 36480
rect 16480 35392 16800 36416
rect 16480 35328 16488 35392
rect 16552 35328 16568 35392
rect 16632 35328 16648 35392
rect 16712 35328 16728 35392
rect 16792 35328 16800 35392
rect 16480 34304 16800 35328
rect 16480 34240 16488 34304
rect 16552 34240 16568 34304
rect 16632 34240 16648 34304
rect 16712 34240 16728 34304
rect 16792 34240 16800 34304
rect 16480 33216 16800 34240
rect 16480 33152 16488 33216
rect 16552 33152 16568 33216
rect 16632 33152 16648 33216
rect 16712 33152 16728 33216
rect 16792 33152 16800 33216
rect 16480 32128 16800 33152
rect 16480 32064 16488 32128
rect 16552 32064 16568 32128
rect 16632 32064 16648 32128
rect 16712 32064 16728 32128
rect 16792 32064 16800 32128
rect 16480 31040 16800 32064
rect 16480 30976 16488 31040
rect 16552 30976 16568 31040
rect 16632 30976 16648 31040
rect 16712 30976 16728 31040
rect 16792 30976 16800 31040
rect 16480 29952 16800 30976
rect 16480 29888 16488 29952
rect 16552 29888 16568 29952
rect 16632 29888 16648 29952
rect 16712 29888 16728 29952
rect 16792 29888 16800 29952
rect 16480 28864 16800 29888
rect 16480 28800 16488 28864
rect 16552 28800 16568 28864
rect 16632 28800 16648 28864
rect 16712 28800 16728 28864
rect 16792 28800 16800 28864
rect 16480 27776 16800 28800
rect 16480 27712 16488 27776
rect 16552 27712 16568 27776
rect 16632 27712 16648 27776
rect 16712 27712 16728 27776
rect 16792 27712 16800 27776
rect 16480 26688 16800 27712
rect 16480 26624 16488 26688
rect 16552 26624 16568 26688
rect 16632 26624 16648 26688
rect 16712 26624 16728 26688
rect 16792 26624 16800 26688
rect 16480 25600 16800 26624
rect 16480 25536 16488 25600
rect 16552 25536 16568 25600
rect 16632 25536 16648 25600
rect 16712 25536 16728 25600
rect 16792 25536 16800 25600
rect 16480 24512 16800 25536
rect 16480 24448 16488 24512
rect 16552 24448 16568 24512
rect 16632 24448 16648 24512
rect 16712 24448 16728 24512
rect 16792 24448 16800 24512
rect 16480 23424 16800 24448
rect 16480 23360 16488 23424
rect 16552 23360 16568 23424
rect 16632 23360 16648 23424
rect 16712 23360 16728 23424
rect 16792 23360 16800 23424
rect 16480 22336 16800 23360
rect 16480 22272 16488 22336
rect 16552 22272 16568 22336
rect 16632 22272 16648 22336
rect 16712 22272 16728 22336
rect 16792 22272 16800 22336
rect 16480 21248 16800 22272
rect 16480 21184 16488 21248
rect 16552 21184 16568 21248
rect 16632 21184 16648 21248
rect 16712 21184 16728 21248
rect 16792 21184 16800 21248
rect 16480 20160 16800 21184
rect 16480 20096 16488 20160
rect 16552 20096 16568 20160
rect 16632 20096 16648 20160
rect 16712 20096 16728 20160
rect 16792 20096 16800 20160
rect 16480 19072 16800 20096
rect 16480 19008 16488 19072
rect 16552 19008 16568 19072
rect 16632 19008 16648 19072
rect 16712 19008 16728 19072
rect 16792 19008 16800 19072
rect 16480 17984 16800 19008
rect 16480 17920 16488 17984
rect 16552 17920 16568 17984
rect 16632 17920 16648 17984
rect 16712 17920 16728 17984
rect 16792 17920 16800 17984
rect 16480 16896 16800 17920
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 16480 14720 16800 15744
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16480 11456 16800 12480
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 16480 10368 16800 11392
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16480 8192 16800 9216
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 7104 16800 8128
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 46816 19019 47376
rect 18699 46752 18707 46816
rect 18771 46752 18787 46816
rect 18851 46752 18867 46816
rect 18931 46752 18947 46816
rect 19011 46752 19019 46816
rect 18699 45728 19019 46752
rect 18699 45664 18707 45728
rect 18771 45664 18787 45728
rect 18851 45664 18867 45728
rect 18931 45664 18947 45728
rect 19011 45664 19019 45728
rect 18699 44640 19019 45664
rect 18699 44576 18707 44640
rect 18771 44576 18787 44640
rect 18851 44576 18867 44640
rect 18931 44576 18947 44640
rect 19011 44576 19019 44640
rect 18699 43552 19019 44576
rect 18699 43488 18707 43552
rect 18771 43488 18787 43552
rect 18851 43488 18867 43552
rect 18931 43488 18947 43552
rect 19011 43488 19019 43552
rect 18699 42464 19019 43488
rect 18699 42400 18707 42464
rect 18771 42400 18787 42464
rect 18851 42400 18867 42464
rect 18931 42400 18947 42464
rect 19011 42400 19019 42464
rect 18699 41376 19019 42400
rect 18699 41312 18707 41376
rect 18771 41312 18787 41376
rect 18851 41312 18867 41376
rect 18931 41312 18947 41376
rect 19011 41312 19019 41376
rect 18699 40288 19019 41312
rect 18699 40224 18707 40288
rect 18771 40224 18787 40288
rect 18851 40224 18867 40288
rect 18931 40224 18947 40288
rect 19011 40224 19019 40288
rect 18699 39200 19019 40224
rect 18699 39136 18707 39200
rect 18771 39136 18787 39200
rect 18851 39136 18867 39200
rect 18931 39136 18947 39200
rect 19011 39136 19019 39200
rect 18699 38112 19019 39136
rect 18699 38048 18707 38112
rect 18771 38048 18787 38112
rect 18851 38048 18867 38112
rect 18931 38048 18947 38112
rect 19011 38048 19019 38112
rect 18699 37024 19019 38048
rect 18699 36960 18707 37024
rect 18771 36960 18787 37024
rect 18851 36960 18867 37024
rect 18931 36960 18947 37024
rect 19011 36960 19019 37024
rect 18699 35936 19019 36960
rect 18699 35872 18707 35936
rect 18771 35872 18787 35936
rect 18851 35872 18867 35936
rect 18931 35872 18947 35936
rect 19011 35872 19019 35936
rect 18699 34848 19019 35872
rect 18699 34784 18707 34848
rect 18771 34784 18787 34848
rect 18851 34784 18867 34848
rect 18931 34784 18947 34848
rect 19011 34784 19019 34848
rect 18699 33760 19019 34784
rect 18699 33696 18707 33760
rect 18771 33696 18787 33760
rect 18851 33696 18867 33760
rect 18931 33696 18947 33760
rect 19011 33696 19019 33760
rect 18699 32672 19019 33696
rect 18699 32608 18707 32672
rect 18771 32608 18787 32672
rect 18851 32608 18867 32672
rect 18931 32608 18947 32672
rect 19011 32608 19019 32672
rect 18699 31584 19019 32608
rect 18699 31520 18707 31584
rect 18771 31520 18787 31584
rect 18851 31520 18867 31584
rect 18931 31520 18947 31584
rect 19011 31520 19019 31584
rect 18699 30496 19019 31520
rect 18699 30432 18707 30496
rect 18771 30432 18787 30496
rect 18851 30432 18867 30496
rect 18931 30432 18947 30496
rect 19011 30432 19019 30496
rect 18699 29408 19019 30432
rect 18699 29344 18707 29408
rect 18771 29344 18787 29408
rect 18851 29344 18867 29408
rect 18931 29344 18947 29408
rect 19011 29344 19019 29408
rect 18699 28320 19019 29344
rect 18699 28256 18707 28320
rect 18771 28256 18787 28320
rect 18851 28256 18867 28320
rect 18931 28256 18947 28320
rect 19011 28256 19019 28320
rect 18699 27232 19019 28256
rect 18699 27168 18707 27232
rect 18771 27168 18787 27232
rect 18851 27168 18867 27232
rect 18931 27168 18947 27232
rect 19011 27168 19019 27232
rect 18699 26144 19019 27168
rect 18699 26080 18707 26144
rect 18771 26080 18787 26144
rect 18851 26080 18867 26144
rect 18931 26080 18947 26144
rect 19011 26080 19019 26144
rect 18699 25056 19019 26080
rect 18699 24992 18707 25056
rect 18771 24992 18787 25056
rect 18851 24992 18867 25056
rect 18931 24992 18947 25056
rect 19011 24992 19019 25056
rect 18699 23968 19019 24992
rect 18699 23904 18707 23968
rect 18771 23904 18787 23968
rect 18851 23904 18867 23968
rect 18931 23904 18947 23968
rect 19011 23904 19019 23968
rect 18699 22880 19019 23904
rect 18699 22816 18707 22880
rect 18771 22816 18787 22880
rect 18851 22816 18867 22880
rect 18931 22816 18947 22880
rect 19011 22816 19019 22880
rect 18699 21792 19019 22816
rect 18699 21728 18707 21792
rect 18771 21728 18787 21792
rect 18851 21728 18867 21792
rect 18931 21728 18947 21792
rect 19011 21728 19019 21792
rect 18699 20704 19019 21728
rect 18699 20640 18707 20704
rect 18771 20640 18787 20704
rect 18851 20640 18867 20704
rect 18931 20640 18947 20704
rect 19011 20640 19019 20704
rect 18699 19616 19019 20640
rect 18699 19552 18707 19616
rect 18771 19552 18787 19616
rect 18851 19552 18867 19616
rect 18931 19552 18947 19616
rect 19011 19552 19019 19616
rect 18699 18528 19019 19552
rect 18699 18464 18707 18528
rect 18771 18464 18787 18528
rect 18851 18464 18867 18528
rect 18931 18464 18947 18528
rect 19011 18464 19019 18528
rect 18699 17440 19019 18464
rect 18699 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19019 17440
rect 18699 16352 19019 17376
rect 18699 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19019 16352
rect 18699 15264 19019 16288
rect 18699 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19019 15264
rect 18699 14176 19019 15200
rect 18699 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19019 14176
rect 18699 13088 19019 14112
rect 18699 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19019 13088
rect 18699 12000 19019 13024
rect 18699 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19019 12000
rect 18699 10912 19019 11936
rect 18699 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19019 10912
rect 18699 9824 19019 10848
rect 18699 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19019 9824
rect 18699 8736 19019 9760
rect 18699 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19019 8736
rect 18699 7648 19019 8672
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1676037725
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_12
timestamp 1676037725
transform 1 0 2208 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_30
timestamp 1676037725
transform 1 0 3864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1676037725
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1676037725
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_48
timestamp 1676037725
transform 1 0 5520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1676037725
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_10
timestamp 1676037725
transform 1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_21
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1676037725
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1676037725
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_78
timestamp 1676037725
transform 1 0 8280 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_90
timestamp 1676037725
transform 1 0 9384 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_102
timestamp 1676037725
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1676037725
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1676037725
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1676037725
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_72
timestamp 1676037725
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_12
timestamp 1676037725
transform 1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1676037725
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_76
timestamp 1676037725
transform 1 0 8096 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_88
timestamp 1676037725
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_100
timestamp 1676037725
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1676037725
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_13
timestamp 1676037725
transform 1 0 2300 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1676037725
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_18
timestamp 1676037725
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_30
timestamp 1676037725
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_76
timestamp 1676037725
transform 1 0 8096 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_88
timestamp 1676037725
transform 1 0 9200 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_100
timestamp 1676037725
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1676037725
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1676037725
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_48
timestamp 1676037725
transform 1 0 5520 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_60
timestamp 1676037725
transform 1 0 6624 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_72
timestamp 1676037725
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_17
timestamp 1676037725
transform 1 0 2668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1676037725
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_76
timestamp 1676037725
transform 1 0 8096 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_88
timestamp 1676037725
transform 1 0 9200 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_100
timestamp 1676037725
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1676037725
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_14
timestamp 1676037725
transform 1 0 2392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_22
timestamp 1676037725
transform 1 0 3128 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp 1676037725
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1676037725
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_10
timestamp 1676037725
transform 1 0 2024 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1676037725
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1676037725
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_13
timestamp 1676037725
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_25
timestamp 1676037725
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_37
timestamp 1676037725
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_78
timestamp 1676037725
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_90
timestamp 1676037725
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_102
timestamp 1676037725
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1676037725
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1676037725
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1676037725
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_71
timestamp 1676037725
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_78
timestamp 1676037725
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_90
timestamp 1676037725
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1676037725
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_70
timestamp 1676037725
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_16
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_23
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1676037725
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_9
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_13
timestamp 1676037725
transform 1 0 2300 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1676037725
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_33
timestamp 1676037725
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_50
timestamp 1676037725
transform 1 0 5704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1676037725
transform 1 0 6440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_75
timestamp 1676037725
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1676037725
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1676037725
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_36
timestamp 1676037725
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1676037725
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_75
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_87
timestamp 1676037725
transform 1 0 9108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_99
timestamp 1676037725
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1676037725
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1676037725
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_26
timestamp 1676037725
transform 1 0 3496 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_34
timestamp 1676037725
transform 1 0 4232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1676037725
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_75
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_87
timestamp 1676037725
transform 1 0 9108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1676037725
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_49
timestamp 1676037725
transform 1 0 5612 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_72
timestamp 1676037725
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1676037725
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1676037725
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_75
timestamp 1676037725
transform 1 0 8004 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_87
timestamp 1676037725
transform 1 0 9108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_99
timestamp 1676037725
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1676037725
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1676037725
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1676037725
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1676037725
transform 1 0 2668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_46
timestamp 1676037725
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_75
timestamp 1676037725
transform 1 0 8004 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_87
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_99
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_8
timestamp 1676037725
transform 1 0 1840 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_16
timestamp 1676037725
transform 1 0 2576 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1676037725
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 1676037725
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1676037725
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1676037725
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_24
timestamp 1676037725
transform 1 0 3312 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_36
timestamp 1676037725
transform 1 0 4416 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_48
timestamp 1676037725
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_189
timestamp 1676037725
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_12
timestamp 1676037725
transform 1 0 2208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_16
timestamp 1676037725
transform 1 0 2576 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_189
timestamp 1676037725
transform 1 0 18492 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1676037725
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_23
timestamp 1676037725
transform 1 0 3220 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1676037725
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_43
timestamp 1676037725
transform 1 0 5060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1676037725
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1676037725
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_7
timestamp 1676037725
transform 1 0 1748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_12
timestamp 1676037725
transform 1 0 2208 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_18
timestamp 1676037725
transform 1 0 2760 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1676037725
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_52
timestamp 1676037725
transform 1 0 5888 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_64
timestamp 1676037725
transform 1 0 6992 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_45
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1676037725
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_65
timestamp 1676037725
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_88
timestamp 1676037725
transform 1 0 9200 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1676037725
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_189
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 1676037725
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_39
timestamp 1676037725
transform 1 0 4692 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_52
timestamp 1676037725
transform 1 0 5888 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_64
timestamp 1676037725
transform 1 0 6992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_68
timestamp 1676037725
transform 1 0 7360 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1676037725
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1676037725
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_70
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1676037725
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_49
timestamp 1676037725
transform 1 0 5612 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_54
timestamp 1676037725
transform 1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_64
timestamp 1676037725
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1676037725
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_189
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1676037725
transform 1 0 1840 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_20
timestamp 1676037725
transform 1 0 2944 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_37
timestamp 1676037725
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1676037725
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_66
timestamp 1676037725
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_75
timestamp 1676037725
transform 1 0 8004 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_87
timestamp 1676037725
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_99
timestamp 1676037725
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_189
timestamp 1676037725
transform 1 0 18492 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1676037725
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_14
timestamp 1676037725
transform 1 0 2392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1676037725
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_52
timestamp 1676037725
transform 1 0 5888 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_60
timestamp 1676037725
transform 1 0 6624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1676037725
transform 1 0 7544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1676037725
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_23
timestamp 1676037725
transform 1 0 3220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_33
timestamp 1676037725
transform 1 0 4140 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_41
timestamp 1676037725
transform 1 0 4876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1676037725
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_65
timestamp 1676037725
transform 1 0 7084 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_71
timestamp 1676037725
transform 1 0 7636 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_77
timestamp 1676037725
transform 1 0 8188 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_89
timestamp 1676037725
transform 1 0 9292 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_101
timestamp 1676037725
transform 1 0 10396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1676037725
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_189
timestamp 1676037725
transform 1 0 18492 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 1676037725
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_14
timestamp 1676037725
transform 1 0 2392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1676037725
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_45
timestamp 1676037725
transform 1 0 5244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_52
timestamp 1676037725
transform 1 0 5888 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_61
timestamp 1676037725
transform 1 0 6716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1676037725
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_34
timestamp 1676037725
transform 1 0 4232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_46
timestamp 1676037725
transform 1 0 5336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1676037725
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_66
timestamp 1676037725
transform 1 0 7176 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_90
timestamp 1676037725
transform 1 0 9384 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_102
timestamp 1676037725
transform 1 0 10488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1676037725
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_189
timestamp 1676037725
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_33
timestamp 1676037725
transform 1 0 4140 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_44
timestamp 1676037725
transform 1 0 5152 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_50
timestamp 1676037725
transform 1 0 5704 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_56
timestamp 1676037725
transform 1 0 6256 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_67
timestamp 1676037725
transform 1 0 7268 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_79
timestamp 1676037725
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1676037725
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1676037725
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_33
timestamp 1676037725
transform 1 0 4140 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_47
timestamp 1676037725
transform 1 0 5428 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1676037725
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_68
timestamp 1676037725
transform 1 0 7360 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_74
timestamp 1676037725
transform 1 0 7912 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_82
timestamp 1676037725
transform 1 0 8648 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_94
timestamp 1676037725
transform 1 0 9752 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 1676037725
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_189
timestamp 1676037725
transform 1 0 18492 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_21
timestamp 1676037725
transform 1 0 3036 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1676037725
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_77
timestamp 1676037725
transform 1 0 8188 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_85
timestamp 1676037725
transform 1 0 8924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_97
timestamp 1676037725
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1676037725
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_189
timestamp 1676037725
transform 1 0 18492 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1676037725
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_33
timestamp 1676037725
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_63
timestamp 1676037725
transform 1 0 6900 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_46
timestamp 1676037725
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1676037725
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_66
timestamp 1676037725
transform 1 0 7176 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_76
timestamp 1676037725
transform 1 0 8096 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_88
timestamp 1676037725
transform 1 0 9200 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_189
timestamp 1676037725
transform 1 0 18492 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_45
timestamp 1676037725
transform 1 0 5244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_64
timestamp 1676037725
transform 1 0 6992 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_71
timestamp 1676037725
transform 1 0 7636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_61
timestamp 1676037725
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_71
timestamp 1676037725
transform 1 0 7636 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_78
timestamp 1676037725
transform 1 0 8280 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_90
timestamp 1676037725
transform 1 0 9384 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_102
timestamp 1676037725
transform 1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_189
timestamp 1676037725
transform 1 0 18492 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1676037725
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1676037725
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_49
timestamp 1676037725
transform 1 0 5612 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_71
timestamp 1676037725
transform 1 0 7636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp 1676037725
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1676037725
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_66
timestamp 1676037725
transform 1 0 7176 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_78
timestamp 1676037725
transform 1 0 8280 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_90
timestamp 1676037725
transform 1 0 9384 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_102
timestamp 1676037725
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1676037725
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_189
timestamp 1676037725
transform 1 0 18492 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_33
timestamp 1676037725
transform 1 0 4140 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_56
timestamp 1676037725
transform 1 0 6256 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_68
timestamp 1676037725
transform 1 0 7360 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1676037725
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_43
timestamp 1676037725
transform 1 0 5060 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1676037725
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_189
timestamp 1676037725
transform 1 0 18492 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_63
timestamp 1676037725
transform 1 0 6900 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_75
timestamp 1676037725
transform 1 0 8004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_189
timestamp 1676037725
transform 1 0 18492 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1676037725
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1676037725
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_64
timestamp 1676037725
transform 1 0 6992 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_73
timestamp 1676037725
transform 1 0 7820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 1676037725
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_74
timestamp 1676037725
transform 1 0 7912 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_86
timestamp 1676037725
transform 1 0 9016 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_98
timestamp 1676037725
transform 1 0 10120 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1676037725
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_189
timestamp 1676037725
transform 1 0 18492 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_49
timestamp 1676037725
transform 1 0 5612 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_68
timestamp 1676037725
transform 1 0 7360 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1676037725
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_35
timestamp 1676037725
transform 1 0 4324 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_41
timestamp 1676037725
transform 1 0 4876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1676037725
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_189
timestamp 1676037725
transform 1 0 18492 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_49
timestamp 1676037725
transform 1 0 5612 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_64
timestamp 1676037725
transform 1 0 6992 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_76
timestamp 1676037725
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_189
timestamp 1676037725
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_8
timestamp 1676037725
transform 1 0 1840 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_20
timestamp 1676037725
transform 1 0 2944 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_32
timestamp 1676037725
transform 1 0 4048 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_44
timestamp 1676037725
transform 1 0 5152 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_189
timestamp 1676037725
transform 1 0 18492 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_189
timestamp 1676037725
transform 1 0 18492 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_189
timestamp 1676037725
transform 1 0 18492 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_9
timestamp 1676037725
transform 1 0 1932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1676037725
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1676037725
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1676037725
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_189
timestamp 1676037725
transform 1 0 18492 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_189
timestamp 1676037725
transform 1 0 18492 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_189
timestamp 1676037725
transform 1 0 18492 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_189
timestamp 1676037725
transform 1 0 18492 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_8
timestamp 1676037725
transform 1 0 1840 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_20
timestamp 1676037725
transform 1 0 2944 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1676037725
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_189
timestamp 1676037725
transform 1 0 18492 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_189
timestamp 1676037725
transform 1 0 18492 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_189
timestamp 1676037725
transform 1 0 18492 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_9
timestamp 1676037725
transform 1 0 1932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1676037725
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_57
timestamp 1676037725
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_69
timestamp 1676037725
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1676037725
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_113
timestamp 1676037725
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_125
timestamp 1676037725
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1676037725
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_169
timestamp 1676037725
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_181
timestamp 1676037725
transform 1 0 17756 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 18860 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 18860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 18860 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 18860 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 18860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 18860 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 18860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _107_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _108_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _109_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _110_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _111_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _112_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _113_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3036 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _114_
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _115_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2392 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _116_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _117_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3128 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _118_
timestamp 1676037725
transform -1 0 2208 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _119_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _120_
timestamp 1676037725
transform 1 0 1840 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _121_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3128 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _122_
timestamp 1676037725
transform -1 0 2760 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _123_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7636 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1676037725
transform 1 0 8096 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1676037725
transform -1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _126_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _127_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7084 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _128_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _129_
timestamp 1676037725
transform 1 0 2852 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _130_
timestamp 1676037725
transform 1 0 2852 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _131_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3496 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _132_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_2  _133_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5152 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or4b_2  _134_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _135_
timestamp 1676037725
transform -1 0 4232 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_2  _136_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and4_4  _137_
timestamp 1676037725
transform -1 0 7360 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _138_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _139_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _140_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7636 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _141_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5888 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1676037725
transform 1 0 8004 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _143_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6900 0 1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_8  _144_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7360 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__a31o_1  _145_
timestamp 1676037725
transform 1 0 6532 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _146_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6992 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_4  _147_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6072 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_2  _148_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8188 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _149_
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_2  _150_
timestamp 1676037725
transform -1 0 8924 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _151_
timestamp 1676037725
transform -1 0 8188 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _152_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _153_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__nand2_2  _154_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4876 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _155_
timestamp 1676037725
transform -1 0 5888 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _156_
timestamp 1676037725
transform -1 0 7176 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _157_
timestamp 1676037725
transform -1 0 7820 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_2  _158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6992 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o311ai_4  _159_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7636 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _160_
timestamp 1676037725
transform 1 0 7544 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _161_
timestamp 1676037725
transform 1 0 6256 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _162_
timestamp 1676037725
transform 1 0 6624 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _163_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7544 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _164_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6256 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_2  _165_
timestamp 1676037725
transform -1 0 8556 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _166_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8004 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _167_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5336 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _168_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8464 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _169_
timestamp 1676037725
transform -1 0 5612 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _170_
timestamp 1676037725
transform 1 0 5336 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1676037725
transform -1 0 4692 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _172_
timestamp 1676037725
transform -1 0 5888 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _173_
timestamp 1676037725
transform 1 0 4140 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _174_
timestamp 1676037725
transform 1 0 3496 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _175_
timestamp 1676037725
transform -1 0 2208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _176_
timestamp 1676037725
transform 1 0 2668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _177_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _178_
timestamp 1676037725
transform -1 0 2392 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _179_
timestamp 1676037725
transform 1 0 2576 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _180_
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _181_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _182_
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _183_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5244 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _184_
timestamp 1676037725
transform -1 0 4876 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _185_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _186_
timestamp 1676037725
transform 1 0 7452 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _187_
timestamp 1676037725
transform -1 0 8372 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp 1676037725
transform -1 0 8004 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _189_
timestamp 1676037725
transform 1 0 5520 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_4  _190_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7176 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_1  _191_
timestamp 1676037725
transform -1 0 6716 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _192_
timestamp 1676037725
transform -1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _193_
timestamp 1676037725
transform 1 0 5796 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _194_
timestamp 1676037725
transform -1 0 6072 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _195_
timestamp 1676037725
transform 1 0 3128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _196_
timestamp 1676037725
transform 1 0 4048 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _197_
timestamp 1676037725
transform -1 0 4140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _198_
timestamp 1676037725
transform 1 0 2760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _199_
timestamp 1676037725
transform 1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _200_
timestamp 1676037725
transform -1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _201_
timestamp 1676037725
transform -1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _202_
timestamp 1676037725
transform 1 0 2392 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _203_
timestamp 1676037725
transform -1 0 3128 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _204_
timestamp 1676037725
transform 1 0 2208 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _205_
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _206_
timestamp 1676037725
transform -1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1676037725
transform 1 0 2760 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _208_
timestamp 1676037725
transform 1 0 2852 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _209_
timestamp 1676037725
transform -1 0 3956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _210_
timestamp 1676037725
transform -1 0 3312 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _211_
timestamp 1676037725
transform -1 0 2300 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _212_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _213_
timestamp 1676037725
transform -1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _214_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6072 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _215_
timestamp 1676037725
transform 1 0 6440 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _216_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1676037725
transform -1 0 5428 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1676037725
transform -1 0 6072 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1676037725
transform -1 0 3496 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _221_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _222_
timestamp 1676037725
transform 1 0 6532 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _223_
timestamp 1676037725
transform 1 0 3772 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _225_
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _226_
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _227_
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _228_
timestamp 1676037725
transform 1 0 3956 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _229_
timestamp 1676037725
transform 1 0 4232 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _230_
timestamp 1676037725
transform -1 0 8096 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _231_
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _232_
timestamp 1676037725
transform 1 0 6164 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _233_
timestamp 1676037725
transform -1 0 5612 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _234_
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1676037725
transform 1 0 6532 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _236_
timestamp 1676037725
transform 1 0 6164 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _237_
timestamp 1676037725
transform 1 0 3772 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1676037725
transform -1 0 3772 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1676037725
transform -1 0 5428 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _240_
timestamp 1676037725
transform -1 0 5888 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _241_
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp 1676037725
transform -1 0 5704 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _243_
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _244_
timestamp 1676037725
transform -1 0 5520 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _245_
timestamp 1676037725
transform -1 0 8280 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _246_
timestamp 1676037725
transform 1 0 6532 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _247_
timestamp 1676037725
transform 1 0 6256 0 1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _248_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 5244 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6440 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7176 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  max_cap11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output3
timestamp 1676037725
transform -1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output4
timestamp 1676037725
transform -1 0 1932 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1676037725
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1676037725
transform -1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1676037725
transform -1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1676037725
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  segment7_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 1840 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  segment7_13
timestamp 1676037725
transform -1 0 1840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  segment7_14
timestamp 1676037725
transform -1 0 1840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  segment7_15
timestamp 1676037725
transform -1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  segment7_16
timestamp 1676037725
transform -1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  segment7_17
timestamp 1676037725
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  segment7_18
timestamp 1676037725
transform -1 0 2576 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 47880 800 48000 0 FreeSans 480 0 0 0 led_out[0]
port 1 nsew signal tristate
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 led_out[1]
port 2 nsew signal tristate
flabel metal3 s 0 33736 800 33856 0 FreeSans 480 0 0 0 led_out[2]
port 3 nsew signal tristate
flabel metal3 s 0 26664 800 26784 0 FreeSans 480 0 0 0 led_out[3]
port 4 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 led_out[4]
port 5 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 led_out[5]
port 6 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 led_out[6]
port 7 nsew signal tristate
flabel metal3 s 0 44344 800 44464 0 FreeSans 480 0 0 0 led_out_b[0]
port 8 nsew signal tristate
flabel metal3 s 0 37272 800 37392 0 FreeSans 480 0 0 0 led_out_b[1]
port 9 nsew signal tristate
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 led_out_b[2]
port 10 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 led_out_b[3]
port 11 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 led_out_b[4]
port 12 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 led_out_b[5]
port 13 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 led_out_b[6]
port 14 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 reset
port 15 nsew signal input
flabel metal4 s 3163 2128 3483 47376 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 7602 2128 7922 47376 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 12041 2128 12361 47376 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 16480 2128 16800 47376 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 5382 2128 5702 47376 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 9821 2128 10141 47376 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 14260 2128 14580 47376 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 18699 2128 19019 47376 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 50000
<< end >>
